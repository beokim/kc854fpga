library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bootrom is
    generic(
        ADDR_WIDTH   : integer := 9
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end bootrom;

architecture rtl of bootrom is
    type rom512x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom512x8 := (
         x"3e",  x"4f",  x"d3",  x"8a",  x"3e",  x"15",  x"d3",  x"88", -- 0000
         x"3e",  x"0f",  x"d3",  x"8a",  x"3e",  x"03",  x"d3",  x"8a", -- 0008
         x"3e",  x"08",  x"d3",  x"84",  x"21",  x"00",  x"80",  x"11", -- 0010
         x"01",  x"80",  x"01",  x"00",  x"08",  x"36",  x"33",  x"ed", -- 0018
         x"b0",  x"01",  x"00",  x"08",  x"36",  x"55",  x"ed",  x"b0", -- 0020
         x"01",  x"00",  x"08",  x"36",  x"00",  x"ed",  x"b0",  x"01", -- 0028
         x"00",  x"08",  x"36",  x"0f",  x"ed",  x"b0",  x"01",  x"00", -- 0030
         x"01",  x"36",  x"00",  x"ed",  x"b0",  x"01",  x"00",  x"01", -- 0038
         x"36",  x"ff",  x"ed",  x"b0",  x"01",  x"00",  x"01",  x"36", -- 0040
         x"00",  x"ed",  x"b0",  x"01",  x"00",  x"01",  x"36",  x"ff", -- 0048
         x"ed",  x"b0",  x"01",  x"00",  x"01",  x"36",  x"00",  x"ed", -- 0050
         x"b0",  x"01",  x"00",  x"01",  x"36",  x"ff",  x"ed",  x"b0", -- 0058
         x"01",  x"00",  x"01",  x"36",  x"00",  x"ed",  x"b0",  x"01", -- 0060
         x"ff",  x"00",  x"36",  x"ff",  x"ed",  x"b0",  x"21",  x"00", -- 0068
         x"80",  x"7c",  x"fe",  x"a8",  x"28",  x"21",  x"7d",  x"e6", -- 0070
         x"c1",  x"fe",  x"00",  x"28",  x"15",  x"7d",  x"e6",  x"c2", -- 0078
         x"fe",  x"40",  x"28",  x"0e",  x"7d",  x"e6",  x"c4",  x"fe", -- 0080
         x"80",  x"28",  x"07",  x"7d",  x"e6",  x"c8",  x"fe",  x"c0", -- 0088
         x"20",  x"02",  x"36",  x"00",  x"23",  x"18",  x"da",  x"21", -- 0090
         x"40",  x"8f",  x"11",  x"c0",  x"00",  x"0e",  x"08",  x"af", -- 0098
         x"06",  x"40",  x"19",  x"77",  x"3c",  x"23",  x"10",  x"fb", -- 00A0
         x"0d",  x"20",  x"f5",  x"21",  x"7f",  x"8f",  x"11",  x"00", -- 00A8
         x"01",  x"0e",  x"08",  x"3e",  x"80",  x"06",  x"08",  x"19", -- 00B0
         x"77",  x"0f",  x"2b",  x"10",  x"fb",  x"0d",  x"20",  x"f5", -- 00B8
         x"21",  x"00",  x"90",  x"cb",  x"5c",  x"20",  x"10",  x"7d", -- 00C0
         x"e6",  x"c0",  x"fe",  x"c0",  x"20",  x"02",  x"36",  x"ff", -- 00C8
         x"23",  x"18",  x"f0",  x"3e",  x"3f",  x"d3",  x"88",  x"3e", -- 00D0
         x"0a",  x"d3",  x"84",  x"21",  x"00",  x"80",  x"11",  x"01", -- 00D8
         x"80",  x"01",  x"ff",  x"27",  x"36",  x"39",  x"ed",  x"b0", -- 00E0
         x"21",  x"00",  x"94",  x"7c",  x"fe",  x"98",  x"28",  x"0c", -- 00E8
         x"7d",  x"e6",  x"c0",  x"fe",  x"00",  x"20",  x"02",  x"36", -- 00F0
         x"99",  x"23",  x"18",  x"ef",  x"21",  x"00",  x"90",  x"11", -- 00F8
         x"80",  x"00",  x"0e",  x"08",  x"af",  x"06",  x"80",  x"19", -- 0100
         x"cb",  x"b7",  x"cb",  x"6d",  x"28",  x"02",  x"cb",  x"f7", -- 0108
         x"77",  x"23",  x"10",  x"f4",  x"c6",  x"09",  x"0d",  x"20", -- 0110
         x"ec",  x"3e",  x"45",  x"d3",  x"8e",  x"3e",  x"19",  x"d3", -- 0118
         x"8e",  x"18",  x"fe",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0120
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0128
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0130
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0138
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0140
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0148
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0150
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0158
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0160
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0168
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0170
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0178
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0180
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0188
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0190
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0198
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 01F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 01F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
