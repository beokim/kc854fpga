library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bootrom is
    generic(
        ADDR_WIDTH   : integer := 10
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end bootrom;

architecture rtl of bootrom is
    type rom1024x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom1024x8 := (
         x"3e",  x"4f",  x"d3",  x"8a",  x"3e",  x"15",  x"d3",  x"88", -- 0000
         x"3e",  x"0f",  x"d3",  x"8a",  x"3e",  x"03",  x"d3",  x"8a", -- 0008
         x"3e",  x"08",  x"d3",  x"84",  x"21",  x"00",  x"80",  x"11", -- 0010
         x"01",  x"80",  x"01",  x"00",  x"28",  x"36",  x"00",  x"ed", -- 0018
         x"b0",  x"31",  x"00",  x"c0",  x"21",  x"85",  x"00",  x"11", -- 0020
         x"00",  x"80",  x"cd",  x"40",  x"00",  x"3e",  x"0a",  x"d3", -- 0028
         x"84",  x"21",  x"00",  x"80",  x"11",  x"01",  x"80",  x"01", -- 0030
         x"ff",  x"27",  x"36",  x"39",  x"ed",  x"b0",  x"18",  x"fe", -- 0038
         x"3e",  x"80",  x"ed",  x"a0",  x"cd",  x"7f",  x"00",  x"30", -- 0040
         x"f9",  x"d5",  x"01",  x"00",  x"00",  x"50",  x"14",  x"cd", -- 0048
         x"7f",  x"00",  x"30",  x"fa",  x"d4",  x"7f",  x"00",  x"cb", -- 0050
         x"11",  x"cb",  x"10",  x"38",  x"1f",  x"15",  x"20",  x"f4", -- 0058
         x"03",  x"5e",  x"23",  x"cb",  x"33",  x"30",  x"0c",  x"16", -- 0060
         x"10",  x"cd",  x"7f",  x"00",  x"cb",  x"12",  x"30",  x"f9", -- 0068
         x"14",  x"cb",  x"3a",  x"cb",  x"1b",  x"e3",  x"e5",  x"ed", -- 0070
         x"52",  x"d1",  x"ed",  x"b0",  x"e1",  x"30",  x"c5",  x"87", -- 0078
         x"c0",  x"7e",  x"23",  x"17",  x"c9",  x"00",  x"9c",  x"00", -- 0080
         x"66",  x"3c",  x"14",  x"ff",  x"3c",  x"66",  x"07",  x"c6", -- 0088
         x"04",  x"cc",  x"18",  x"30",  x"66",  x"c6",  x"04",  x"8c", -- 0090
         x"07",  x"0c",  x"c1",  x"00",  x"fc",  x"66",  x"66",  x"7c", -- 0098
         x"a4",  x"02",  x"fc",  x"07",  x"00",  x"6c",  x"66",  x"e6", -- 00A0
         x"00",  x"7c",  x"c6",  x"f0",  x"3c",  x"03",  x"0e",  x"c6", -- 00A8
         x"7c",  x"00",  x"1e",  x"0c",  x"00",  x"18",  x"cc",  x"cc", -- 00B0
         x"78",  x"8e",  x"07",  x"ee",  x"fe",  x"d6",  x"c6",  x"00", -- 00B8
         x"11",  x"17",  x"e0",  x"13",  x"14",  x"78",  x"30",  x"30", -- 00C0
         x"00",  x"f0",  x"61",  x"60",  x"00",  x"62",  x"66",  x"fe", -- 00C8
         x"00",  x"8b",  x"c3",  x"c0",  x"00",  x"c4",  x"cb",  x"00", -- 00D0
         x"f8",  x"f2",  x"3c",  x"00",  x"6c",  x"f8",  x"22",  x"2f", -- 00D8
         x"86",  x"03",  x"d6",  x"fe",  x"ee",  x"07",  x"e6",  x"d7", -- 00E0
         x"14",  x"70",  x"57",  x"3c",  x"07",  x"2f",  x"4f",  x"3c", -- 00E8
         x"07",  x"a8",  x"00",  x"7f",  x"18",  x"02",  x"f7",  x"70", -- 00F0
         x"8f",  x"36",  x"30",  x"78",  x"78",  x"fc",  x"02",  x"00", -- 00F8
         x"01",  x"fe",  x"62",  x"68",  x"78",  x"68",  x"62",  x"fe", -- 0100
         x"38",  x"b7",  x"58",  x"8f",  x"58",  x"92",  x"44",  x"47", -- 0108
         x"17",  x"94",  x"27",  x"38",  x"6c",  x"29",  x"6c",  x"44", -- 0110
         x"38",  x"61",  x"07",  x"bb",  x"7c",  x"00",  x"2f",  x"7c", -- 0118
         x"0f",  x"f1",  x"2f",  x"f7",  x"37",  x"5c",  x"78",  x"1f", -- 0120
         x"56",  x"0c",  x"38",  x"60",  x"e2",  x"59",  x"20",  x"07", -- 0128
         x"67",  x"00",  x"9c",  x"b7",  x"a7",  x"87",  x"29",  x"ce", -- 0130
         x"87",  x"70",  x"b7",  x"88",  x"c7",  x"20",  x"e6",  x"f6", -- 0138
         x"de",  x"ce",  x"a9",  x"07",  x"ca",  x"9f",  x"e2",  x"27", -- 0140
         x"c6",  x"b7",  x"73",  x"87",  x"9e",  x"47",  x"73",  x"87", -- 0148
         x"8b",  x"37",  x"b9",  x"4f",  x"e7",  x"07",  x"1f",  x"9c", -- 0150
         x"2f",  x"1c",  x"3c",  x"04",  x"6c",  x"cc",  x"fe",  x"0c", -- 0158
         x"1e",  x"44",  x"07",  x"0d",  x"4b",  x"00",  x"fe",  x"04", -- 0160
         x"9c",  x"ef",  x"27",  x"cf",  x"02",  x"fc",  x"b4",  x"5b", -- 0168
         x"0f",  x"e7",  x"0c",  x"d9",  x"11",  x"f0",  x"e7",  x"87", -- 0170
         x"3c",  x"2f",  x"e1",  x"c7",  x"39",  x"cf",  x"4f",  x"2f", -- 0178
         x"1f",  x"1f",  x"3c",  x"6b",  x"e3",  x"a7",  x"3c",  x"4f", -- 0180
         x"f3",  x"67",  x"cf",  x"3f",  x"2f",  x"03",  x"81",  x"ff", -- 0188
         x"47",  x"9c",  x"87",  x"f0",  x"0f",  x"bc",  x"00",  x"83", -- 0190
         x"87",  x"84",  x"e7",  x"f3",  x"0e",  x"9c",  x"8f",  x"e1", -- 0198
         x"df",  x"3c",  x"1f",  x"e1",  x"d7",  x"3c",  x"26",  x"e3", -- 01A0
         x"97",  x"1a",  x"27",  x"62",  x"89",  x"8f",  x"19",  x"e0", -- 01A8
         x"07",  x"67",  x"00",  x"9c",  x"ef",  x"a3",  x"c3",  x"9f", -- 01B0
         x"12",  x"b4",  x"16",  x"cc",  x"31",  x"37",  x"3a",  x"c7", -- 01B8
         x"42",  x"f3",  x"4f",  x"ce",  x"1f",  x"c7",  x"f3",  x"ce", -- 01C0
         x"00",  x"df",  x"33",  x"ce",  x"00",  x"df",  x"b1",  x"e7", -- 01C8
         x"ef",  x"03",  x"3c",  x"00",  x"79",  x"9f",  x"4e",  x"f7", -- 01D0
         x"50",  x"6f",  x"00",  x"0b",  x"8c",  x"97",  x"f3",  x"00", -- 01D8
         x"84",  x"e7",  x"04",  x"3c",  x"00",  x"e5",  x"8f",  x"00", -- 01E0
         x"fb",  x"cf",  x"00",  x"ef",  x"70",  x"1f",  x"95",  x"00", -- 01E8
         x"cf",  x"d0",  x"1e",  x"fd",  x"00",  x"ae",  x"0e",  x"0c", -- 01F0
         x"38",  x"60",  x"b1",  x"90",  x"00",  x"0f",  x"c7",  x"00", -- 01F8
         x"eb",  x"8f",  x"ff",  x"f3",  x"10",  x"00",  x"00",  x"cf", -- 0200
         x"84",  x"00",  x"00",  x"02",  x"00",  x"00",  x"00",  x"00", -- 0208
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0210
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0218
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0220
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0228
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0230
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0238
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0240
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0248
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0250
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0258
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0260
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0268
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0270
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0278
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0280
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0288
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0290
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0298
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 02F8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0300
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0308
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0310
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0318
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0320
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0328
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0330
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0338
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0340
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0348
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0350
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0358
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0360
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0368
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0370
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0378
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0380
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0388
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0390
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 0398
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03A8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03B8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03C0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03C8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03D0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03D8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03E0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03E8
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 03F0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 03F8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
