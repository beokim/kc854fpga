library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bootrom is
    generic(
        ADDR_WIDTH   : integer := 14
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end bootrom;

architecture rtl of bootrom is
    type rom16384x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(7 downto 0); 
    constant romData : rom16384x8 := (
         x"31",  x"00",  x"c0",  x"3e",  x"1f",  x"d3",  x"88",  x"3e", -- 0000
         x"0f",  x"d3",  x"8a",  x"3e",  x"08",  x"d3",  x"84",  x"3e", -- 0008
         x"80",  x"d3",  x"86",  x"21",  x"4a",  x"1c",  x"11",  x"00", -- 0010
         x"c0",  x"cd",  x"38",  x"00",  x"21",  x"55",  x"25",  x"11", -- 0018
         x"00",  x"e0",  x"cd",  x"38",  x"00",  x"af",  x"d3",  x"86", -- 0020
         x"3e",  x"9f",  x"d3",  x"88",  x"21",  x"7d",  x"00",  x"11", -- 0028
         x"00",  x"c0",  x"cd",  x"38",  x"00",  x"c3",  x"00",  x"f0", -- 0030
         x"3e",  x"80",  x"ed",  x"a0",  x"cd",  x"77",  x"00",  x"30", -- 0038
         x"f9",  x"d5",  x"01",  x"00",  x"00",  x"50",  x"14",  x"cd", -- 0040
         x"77",  x"00",  x"30",  x"fa",  x"d4",  x"77",  x"00",  x"cb", -- 0048
         x"11",  x"cb",  x"10",  x"38",  x"1f",  x"15",  x"20",  x"f4", -- 0050
         x"03",  x"5e",  x"23",  x"cb",  x"33",  x"30",  x"0c",  x"16", -- 0058
         x"10",  x"cd",  x"77",  x"00",  x"cb",  x"12",  x"30",  x"f9", -- 0060
         x"14",  x"cb",  x"3a",  x"cb",  x"1b",  x"e3",  x"e5",  x"ed", -- 0068
         x"52",  x"d1",  x"ed",  x"b0",  x"e1",  x"30",  x"c5",  x"87", -- 0070
         x"c0",  x"7e",  x"23",  x"17",  x"c9",  x"18",  x"00",  x"0b", -- 0078
         x"c3",  x"8c",  x"c0",  x"7f",  x"7f",  x"42",  x"41",  x"00", -- 0080
         x"53",  x"49",  x"43",  x"00",  x"21",  x"bd",  x"c0",  x"11", -- 0088
         x"00",  x"00",  x"03",  x"01",  x"67",  x"00",  x"ed",  x"b0", -- 0090
         x"eb",  x"00",  x"f9",  x"cd",  x"69",  x"c6",  x"32",  x"ab", -- 0098
         x"03",  x"32",  x"00",  x"00",  x"04",  x"21",  x"92",  x"c0", -- 00A0
         x"cd",  x"c9",  x"d1",  x"2c",  x"21",  x"ae",  x"05",  x"cd", -- 00A8
         x"ae",  x"00",  x"c5",  x"21",  x"62",  x"03",  x"cd",  x"86", -- 00B0
         x"c9",  x"7a",  x"18",  x"d6",  x"06",  x"21",  x"2a",  x"2b", -- 00B8
         x"30",  x"03",  x"00",  x"11",  x"ff",  x"bf",  x"23",  x"cd", -- 00C0
         x"89",  x"c6",  x"28",  x"00",  x"09",  x"7e",  x"47",  x"2f", -- 00C8
         x"77",  x"be",  x"70",  x"28",  x"30",  x"f2",  x"2b",  x"42", -- 00D0
         x"ff",  x"22",  x"b0",  x"03",  x"18",  x"19",  x"22",  x"56", -- 00D8
         x"27",  x"41",  x"c6",  x"2a",  x"c0",  x"05",  x"11",  x"ef", -- 00E0
         x"fb",  x"19",  x"cd",  x"29",  x"16",  x"d8",  x"21",  x"a0", -- 00E8
         x"40",  x"2a",  x"00",  x"04",  x"e0",  x"7e",  x"fe",  x"78", -- 00F0
         x"20",  x"01",  x"3e",  x"00",  x"af",  x"32",  x"fc",  x"03", -- 00F8
         x"31",  x"67",  x"03",  x"18",  x"64",  x"0a",  x"7c",  x"52", -- 0100
         x"45",  x"b4",  x"7e",  x"71",  x"c3",  x"00",  x"88",  x"c3", -- 0108
         x"0c",  x"0a",  x"0d",  x"48",  x"43",  x"2d",  x"93",  x"11", -- 0110
         x"09",  x"00",  x"00",  x"20",  x"42",  x"59",  x"54",  x"45", -- 0118
         x"53",  x"20",  x"6a",  x"46",  x"23",  x"45",  x"0d",  x"00", -- 0120
         x"4d",  x"45",  x"4d",  x"4f",  x"52",  x"59",  x"20",  x"45", -- 0128
         x"00",  x"4e",  x"44",  x"20",  x"3f",  x"20",  x"3a",  x"00", -- 0130
         x"c3",  x"02",  x"89",  x"c0",  x"c3",  x"67",  x"c9",  x"00", -- 0138
         x"c0",  x"00",  x"d6",  x"00",  x"6f",  x"7c",  x"de",  x"00", -- 0140
         x"31",  x"67",  x"78",  x"03",  x"47",  x"3e",  x"00",  x"60", -- 0148
         x"12",  x"35",  x"4a",  x"ca",  x"99",  x"39",  x"00",  x"1c", -- 0150
         x"76",  x"98",  x"22",  x"95",  x"b3",  x"98",  x"0a",  x"00", -- 0158
         x"dd",  x"47",  x"98",  x"53",  x"d1",  x"99",  x"99",  x"0a", -- 0160
         x"00",  x"1a",  x"9f",  x"98",  x"65",  x"bc",  x"cd",  x"98", -- 0168
         x"d6",  x"00",  x"77",  x"3e",  x"98",  x"52",  x"c7",  x"4f", -- 0170
         x"80",  x"0b",  x"0f",  x"ff",  x"1b",  x"00",  x"0a",  x"01", -- 0178
         x"2c",  x"f0",  x"49",  x"d7",  x"4e",  x"00",  x"00",  x"65", -- 0180
         x"0b",  x"04",  x"fe",  x"ff",  x"00",  x"43",  x"29",  x"01", -- 0188
         x"04",  x"0d",  x"c5",  x"b0",  x"6b",  x"c6",  x"73",  x"ce", -- 0190
         x"45",  x"58",  x"54",  x"00",  x"c4",  x"41",  x"54",  x"41", -- 0198
         x"c9",  x"4e",  x"50",  x"55",  x"c0",  x"08",  x"49",  x"4d", -- 01A0
         x"d2",  x"45",  x"41",  x"44",  x"18",  x"cc",  x"45",  x"54", -- 01A8
         x"43",  x"54",  x"4f",  x"d2",  x"0d",  x"55",  x"4e",  x"c9", -- 01B0
         x"46",  x"0f",  x"53",  x"e1",  x"09",  x"a3",  x"8c",  x"0f", -- 01B8
         x"53",  x"55",  x"42",  x"0b",  x"54",  x"55",  x"33",  x"52", -- 01C0
         x"4e",  x"05",  x"4d",  x"d3",  x"12",  x"30",  x"50",  x"cf", -- 01C8
         x"2e",  x"cf",  x"4e",  x"ce",  x"55",  x"06",  x"4c",  x"4c", -- 01D0
         x"d7",  x"41",  x"49",  x"38",  x"45",  x"02",  x"46",  x"d0", -- 01D8
         x"4f",  x"4b",  x"45",  x"c4",  x"98",  x"03",  x"c1",  x"17", -- 01E0
         x"4f",  x"cc",  x"49",  x"60",  x"4e",  x"36",  x"c3",  x"4c", -- 01E8
         x"53",  x"d7",  x"49",  x"00",  x"44",  x"54",  x"48",  x"c2", -- 01F0
         x"59",  x"45",  x"a1",  x"c3",  x"66",  x"41",  x"27",  x"d0", -- 01F8
         x"52",  x"15",  x"54",  x"3f",  x"c3",  x"4f",  x"03",  x"1d", -- 0200
         x"52",  x"f6",  x"1c",  x"67",  x"52",  x"04",  x"4f",  x"c1", -- 0208
         x"6c",  x"c3",  x"53",  x"41",  x"56",  x"45",  x"80",  x"85", -- 0210
         x"57",  x"d4",  x"41",  x"00",  x"42",  x"28",  x"d4",  x"4f", -- 0218
         x"c6",  x"4e",  x"d3",  x"50",  x"67",  x"43",  x"07",  x"48", -- 0220
         x"45",  x"5a",  x"86",  x"81",  x"66",  x"45",  x"01",  x"50", -- 0228
         x"ab",  x"ad",  x"aa",  x"af",  x"de",  x"c1",  x"80",  x"aa", -- 0230
         x"cf",  x"52",  x"be",  x"0c",  x"bd",  x"bc",  x"d3",  x"47", -- 0238
         x"91",  x"30",  x"3f",  x"c1",  x"42",  x"53",  x"d5",  x"18", -- 0240
         x"53",  x"52",  x"c6",  x"94",  x"50",  x"b3",  x"60",  x"75", -- 0248
         x"53",  x"d3",  x"51",  x"52",  x"d2",  x"c1",  x"1f",  x"cc", -- 0250
         x"4e",  x"c5",  x"58",  x"50",  x"fe",  x"5d",  x"0d",  x"64", -- 0258
         x"49",  x"4e",  x"0c",  x"c1",  x"54",  x"4e",  x"d0",  x"d7", -- 0260
         x"4a",  x"4b",  x"c4",  x"03",  x"1e",  x"d0",  x"49",  x"cc", -- 0268
         x"4c",  x"49",  x"52",  x"30",  x"24",  x"d6",  x"83",  x"07", -- 0270
         x"c1",  x"53",  x"43",  x"c3",  x"48",  x"09",  x"80",  x"10", -- 0278
         x"46",  x"54",  x"24",  x"d2",  x"49",  x"47",  x"48",  x"d8", -- 0280
         x"05",  x"cd",  x"a1",  x"74",  x"0e",  x"85",  x"06",  x"d4", -- 0288
         x"52",  x"98",  x"14",  x"03",  x"46",  x"18",  x"46",  x"c5", -- 0290
         x"44",  x"cd",  x"30",  x"c5",  x"b9",  x"00",  x"45",  x"80", -- 0298
         x"1a",  x"c9",  x"de",  x"c7",  x"dc",  x"cc",  x"00",  x"48", -- 02A0
         x"ca",  x"ec",  x"cb",  x"01",  x"cf",  x"1f",  x"cc",  x"00", -- 02A8
         x"5d",  x"ca",  x"07",  x"ca",  x"eb",  x"c9",  x"cf",  x"ca", -- 02B0
         x"03",  x"df",  x"c8",  x"f6",  x"c9",  x"25",  x"ca",  x"81", -- 02B8
         x"20",  x"18",  x"c9",  x"ec",  x"d3",  x"00",  x"b3",  x"ca", -- 02C0
         x"c0",  x"cb",  x"f7",  x"d3",  x"c4",  x"d0",  x"30",  x"37", -- 02C8
         x"d4",  x"3a",  x"fa",  x"c5",  x"ea",  x"c6",  x"03",  x"d0", -- 02D0
         x"dd",  x"b9",  x"cb",  x"f4",  x"df",  x"1b",  x"00",  x"38", -- 02D8
         x"db",  x"fa",  x"ca",  x"48",  x"c9",  x"f2",  x"c6",  x"00", -- 02E0
         x"aa",  x"c9",  x"43",  x"dc",  x"41",  x"dd",  x"40",  x"c6", -- 02E8
         x"00",  x"2d",  x"c6",  x"b7",  x"c7",  x"b8",  x"c7",  x"e7", -- 02F0
         x"c3",  x"c0",  x"19",  x"a6",  x"d6",  x"70",  x"d7",  x"bc", -- 02F8
         x"d6",  x"00",  x"03",  x"03",  x"90",  x"d0",  x"e3",  x"d3", -- 0300
         x"bd",  x"d0",  x"00",  x"1f",  x"d9",  x"fd",  x"d9",  x"59", -- 0308
         x"d5",  x"6d",  x"d9",  x"00",  x"70",  x"da",  x"76",  x"da", -- 0310
         x"d7",  x"da",  x"ec",  x"da",  x"30",  x"31",  x"d4",  x"86", -- 0318
         x"00",  x"d5",  x"d6",  x"2c",  x"d3",  x"56",  x"d1",  x"bf", -- 0320
         x"d3",  x"00",  x"3b",  x"d3",  x"4b",  x"d3",  x"5b",  x"d3", -- 0328
         x"89",  x"d3",  x"00",  x"92",  x"d3",  x"79",  x"11",  x"d8", -- 0330
         x"79",  x"6a",  x"d4",  x"00",  x"7c",  x"98",  x"d5",  x"7c", -- 0338
         x"f3",  x"d5",  x"7f",  x"28",  x"00",  x"d9",  x"50",  x"5e", -- 0340
         x"ce",  x"46",  x"5d",  x"ce",  x"4e",  x"00",  x"46",  x"53", -- 0348
         x"4e",  x"52",  x"47",  x"4f",  x"44",  x"46",  x"06",  x"43", -- 0350
         x"4f",  x"56",  x"4f",  x"4d",  x"84",  x"58",  x"91",  x"85", -- 0358
         x"44",  x"44",  x"2f",  x"30",  x"0e",  x"ed",  x"c5",  x"6c", -- 0360
         x"53",  x"bc",  x"31",  x"de",  x"0c",  x"43",  x"4e",  x"55", -- 0368
         x"46",  x"0a",  x"49",  x"4f",  x"cd",  x"d0",  x"52",  x"81", -- 0370
         x"d4",  x"52",  x"07",  x"9e",  x"ec",  x"95",  x"21",  x"20", -- 0378
         x"00",  x"46",  x"49",  x"8e",  x"f4",  x"ef",  x"6c",  x"4f", -- 0380
         x"d5",  x"8c",  x"44",  x"0d",  x"a7",  x"b3",  x"f2",  x"62", -- 0388
         x"42",  x"c0",  x"41",  x"00",  x"4b",  x"00",  x"e5",  x"2a", -- 0390
         x"db",  x"03",  x"06",  x"00",  x"00",  x"09",  x"09",  x"3e", -- 0398
         x"e5",  x"3e",  x"d0",  x"95",  x"6f",  x"00",  x"3e",  x"ff", -- 03A0
         x"9c",  x"38",  x"04",  x"67",  x"39",  x"e1",  x"00",  x"d8", -- 03A8
         x"1e",  x"0c",  x"18",  x"14",  x"2a",  x"ca",  x"03",  x"00", -- 03B0
         x"22",  x"58",  x"03",  x"1e",  x"02",  x"01",  x"1e",  x"14", -- 03B8
         x"db",  x"02",  x"00",  x"02",  x"12",  x"02",  x"5a",  x"22", -- 03C0
         x"bb",  x"b4",  x"43",  x"fe",  x"00",  x"55",  x"cb",  x"21", -- 03C8
         x"dd",  x"c2",  x"57",  x"19",  x"44",  x"06",  x"4d",  x"0b", -- 03D0
         x"3e",  x"3f",  x"1e",  x"0e",  x"d6",  x"d4",  x"c4",  x"05", -- 03D8
         x"c3",  x"b5",  x"83",  x"d9",  x"2e",  x"11",  x"e2",  x"d2", -- 03E0
         x"b4",  x"80",  x"ca",  x"0d",  x"c0",  x"7c",  x"a5",  x"3c", -- 03E8
         x"c4",  x"04",  x"21",  x"d8",  x"3e",  x"c1",  x"af",  x"cb", -- 03F0
         x"2f",  x"1d",  x"20",  x"00",  x"37",  x"dc",  x"fd",  x"dd", -- 03F8
         x"cd",  x"df",  x"c6",  x"2b",  x"a0",  x"57",  x"21",  x"ea", -- 0400
         x"03",  x"3a",  x"00",  x"4d",  x"03",  x"b7",  x"28",  x"6b", -- 0408
         x"ed",  x"5b",  x"4e",  x"00",  x"03",  x"f2",  x"f0",  x"c3", -- 0410
         x"d5",  x"cd",  x"2a",  x"d8",  x"60",  x"d1",  x"04",  x"bb", -- 0418
         x"c4",  x"3e",  x"2a",  x"38",  x"1b",  x"02",  x"3e",  x"20", -- 0420
         x"8f",  x"29",  x"c6",  x"92",  x"87",  x"d1",  x"30",  x"06", -- 0428
         x"3f",  x"86",  x"25",  x"18",  x"ba",  x"2a",  x"50",  x"f7", -- 0430
         x"a0",  x"38",  x"f4",  x"d5",  x"11",  x"f9",  x"bc",  x"5d", -- 0438
         x"15",  x"ea",  x"22",  x"e9",  x"33",  x"ae",  x"80",  x"f5", -- 0440
         x"18",  x"47",  x"c8",  x"cd",  x"97",  x"f6",  x"28",  x"b5", -- 0448
         x"28",  x"c0",  x"c1",  x"39",  x"30",  x"58",  x"03",  x"d5", -- 0450
         x"7e",  x"23",  x"b6",  x"23",  x"28",  x"3e",  x"56",  x"7f", -- 0458
         x"34",  x"0a",  x"66",  x"56",  x"6f",  x"26",  x"94",  x"a0", -- 0460
         x"de",  x"d1",  x"c2",  x"96",  x"c3",  x"01",  x"38",  x"b7", -- 0468
         x"3f",  x"18",  x"cd",  x"3e",  x"3e",  x"2b",  x"56",  x"da", -- 0470
         x"0f",  x"30",  x"21",  x"61",  x"19",  x"bd",  x"c8",  x"3c", -- 0478
         x"3d",  x"6a",  x"ca",  x"0a",  x"f5",  x"3f",  x"c0",  x"78", -- 0480
         x"da",  x"c4",  x"47",  x"d1",  x"f1",  x"d2",  x"0d",  x"8a", -- 0488
         x"c8",  x"d5",  x"c5",  x"71",  x"cd",  x"6f",  x"1b",  x"b7", -- 0490
         x"17",  x"52",  x"00",  x"38",  x"08",  x"f1",  x"f5",  x"b7", -- 0498
         x"20",  x"03",  x"c3",  x"00",  x"20",  x"ca",  x"c5",  x"30", -- 04A0
         x"11",  x"eb",  x"2a",  x"d7",  x"05",  x"03",  x"1a",  x"02", -- 04A8
         x"03",  x"13",  x"00",  x"82",  x"20",  x"f7",  x"ed",  x"79", -- 04B0
         x"43",  x"0c",  x"30",  x"28",  x"22",  x"40",  x"13",  x"e3", -- 04B8
         x"c1",  x"09",  x"e5",  x"cd",  x"0c",  x"ab",  x"c4",  x"e1", -- 04C0
         x"22",  x"0a",  x"eb",  x"36",  x"00",  x"ff",  x"d1",  x"23", -- 04C8
         x"23",  x"73",  x"23",  x"72",  x"23",  x"31",  x"11",  x"62", -- 04D0
         x"2b",  x"77",  x"23",  x"13",  x"ef",  x"3c",  x"ef",  x"a0", -- 04D8
         x"d5",  x"23",  x"eb",  x"21",  x"c5",  x"67",  x"e5",  x"62", -- 04E0
         x"6b",  x"01",  x"9e",  x"c8",  x"23",  x"98",  x"04",  x"a6", -- 04E8
         x"3c",  x"05",  x"af",  x"be",  x"23",  x"14",  x"20",  x"fc", -- 04F0
         x"eb",  x"29",  x"18",  x"07",  x"e8",  x"cd",  x"30",  x"c3", -- 04F8
         x"c5",  x"43",  x"40",  x"55",  x"7e",  x"02",  x"c8",  x"0b", -- 0500
         x"2b",  x"06",  x"18",  x"f6",  x"2a",  x"5f",  x"03",  x"d9", -- 0508
         x"34",  x"2a",  x"2b",  x"d6",  x"25",  x"23",  x"c5",  x"14", -- 0510
         x"19",  x"60",  x"58",  x"69",  x"08",  x"3f",  x"c8",  x"3f", -- 0518
         x"18",  x"d0",  x"18",  x"e4",  x"9f",  x"05",  x"af",  x"03", -- 0520
         x"0e",  x"05",  x"6c",  x"5f",  x"08",  x"fb",  x"e5",  x"18", -- 0528
         x"fe",  x"9a",  x"00",  x"71",  x"c5",  x"47",  x"fe",  x"22", -- 0530
         x"ca",  x"91",  x"03",  x"c5",  x"b7",  x"ca",  x"97",  x"c5", -- 0538
         x"3a",  x"1b",  x"00",  x"b7",  x"7e",  x"20",  x"73",  x"fe", -- 0540
         x"3f",  x"3e",  x"9e",  x"36",  x"28",  x"6d",  x"1c",  x"30", -- 0548
         x"ce",  x"41",  x"fe",  x"3c",  x"38",  x"64",  x"88",  x"b8", -- 0550
         x"20",  x"c1",  x"c5",  x"03",  x"01",  x"6d",  x"c5",  x"c5", -- 0558
         x"06",  x"7f",  x"13",  x"07",  x"61",  x"38",  x"07",  x"fe", -- 0560
         x"7b",  x"df",  x"00",  x"e6",  x"5f",  x"77",  x"4e",  x"eb", -- 0568
         x"c0",  x"64",  x"f2",  x"26",  x"c5",  x"04",  x"7e",  x"e6", -- 0570
         x"0e",  x"7f",  x"20",  x"15",  x"3a",  x"b6",  x"06",  x"a7", -- 0578
         x"c8",  x"3a",  x"51",  x"a7",  x"28",  x"c0",  x"3c",  x"57", -- 0580
         x"2a",  x"0c",  x"50",  x"e0",  x"15",  x"c8",  x"b9",  x"20", -- 0588
         x"00",  x"dd",  x"eb",  x"e5",  x"13",  x"1a",  x"b7",  x"fa", -- 0590
         x"69",  x"01",  x"c5",  x"4f",  x"78",  x"fe",  x"88",  x"20", -- 0598
         x"04",  x"42",  x"98",  x"2b",  x"5b",  x"23",  x"43",  x"02", -- 05A0
         x"3f",  x"00",  x"b9",  x"28",  x"e5",  x"e1",  x"18",  x"bb", -- 05A8
         x"48",  x"f1",  x"d4",  x"98",  x"eb",  x"79",  x"60",  x"c1", -- 05B0
         x"f6",  x"12",  x"06",  x"13",  x"0c",  x"d6",  x"3a",  x"28", -- 05B8
         x"6f",  x"49",  x"c6",  x"af",  x"80",  x"a1",  x"d6",  x"54", -- 05C0
         x"03",  x"28",  x"05",  x"d6",  x"0e",  x"c2",  x"e3",  x"d6", -- 05C8
         x"16",  x"7e",  x"e4",  x"41",  x"09",  x"b8",  x"28",  x"e0", -- 05D0
         x"85",  x"1f",  x"0c",  x"13",  x"18",  x"f3",  x"0f",  x"f7", -- 05D8
         x"27",  x"45",  x"01",  x"c9",  x"4c",  x"39",  x"85",  x"00", -- 05E0
         x"52",  x"a1",  x"8c",  x"00",  x"43",  x"4f",  x"92",  x"a5", -- 05E8
         x"86",  x"10",  x"cd",  x"e3",  x"cd",  x"e4",  x"00",  x"dd", -- 05F0
         x"e3",  x"fe",  x"1c",  x"11",  x"9f",  x"c5",  x"28",  x"07", -- 05F8
         x"0e",  x"fe",  x"1d",  x"11",  x"a4",  x"06",  x"80",  x"a7", -- 0600
         x"1e",  x"11",  x"a8",  x"15",  x"c5",  x"20",  x"14",  x"34", -- 0608
         x"8e",  x"c9",  x"cd",  x"2c",  x"a7",  x"cb",  x"6e",  x"a3", -- 0610
         x"80",  x"f1",  x"c5",  x"e1",  x"c3",  x"5e",  x"cb",  x"00", -- 0618
         x"cd",  x"0f",  x"df",  x"20",  x"02",  x"e1",  x"c9",  x"cd", -- 0620
         x"18",  x"27",  x"df",  x"38",  x"e1",  x"87",  x"32",  x"df", -- 0628
         x"18",  x"c1",  x"66",  x"98",  x"8b",  x"d5",  x"dd",  x"23", -- 0630
         x"1c",  x"18",  x"f7",  x"11",  x"f7",  x"0a",  x"d5",  x"28", -- 0638
         x"17",  x"d4",  x"21",  x"eb",  x"e3",  x"28",  x"96",  x"b3", -- 0640
         x"9c",  x"8c",  x"c8",  x"e1",  x"f3",  x"bd",  x"28",  x"28", -- 0648
         x"06",  x"10",  x"c2",  x"48",  x"07",  x"c3",  x"eb",  x"7d", -- 0650
         x"b4",  x"ca",  x"d9",  x"2c",  x"22",  x"10",  x"cb",  x"ff", -- 0658
         x"a3",  x"a3",  x"51",  x"e1",  x"a0",  x"99",  x"c1",  x"c3", -- 0660
         x"9a",  x"03",  x"cd",  x"5f",  x"de",  x"3a",  x"09",  x"91", -- 0668
         x"1c",  x"25",  x"f3",  x"3e",  x"cc",  x"89",  x"b2",  x"dc", -- 0670
         x"05",  x"f1",  x"af",  x"18",  x"ea",  x"c0",  x"16",  x"85", -- 0678
         x"e0",  x"26",  x"5e",  x"03",  x"c3",  x"5d",  x"01",  x"15", -- 0680
         x"d8",  x"68",  x"0d",  x"b5",  x"cf",  x"fa",  x"06",  x"ff", -- 0688
         x"3d",  x"22",  x"c4",  x"17",  x"c3",  x"19",  x"c8",  x"f7", -- 0690
         x"6d",  x"09",  x"d9",  x"02",  x"db",  x"d5",  x"3f",  x"89", -- 0698
         x"e0",  x"97",  x"b4",  x"d8",  x"0a",  x"b2",  x"9a",  x"00", -- 06A0
         x"1d",  x"de",  x"af",  x"6f",  x"67",  x"22",  x"d5",  x"c1", -- 06A8
         x"ff",  x"cc",  x"83",  x"0e",  x"df",  x"03",  x"e5",  x"c5", -- 06B0
         x"2a",  x"31",  x"3b",  x"c9",  x"7c",  x"e5",  x"18",  x"7d", -- 06B8
         x"93",  x"c9",  x"b2",  x"80",  x"41",  x"d8",  x"fe",  x"5b", -- 06C0
         x"3f",  x"c9",  x"3a",  x"f1",  x"51",  x"e5",  x"bb",  x"8f", -- 06C8
         x"79",  x"6e",  x"74",  x"d6",  x"0a",  x"3e",  x"08",  x"18", -- 06D0
         x"eb",  x"4d",  x"fb",  x"0c",  x"dd",  x"f5",  x"de",  x"72", -- 06D8
         x"c8",  x"00",  x"38",  x"13",  x"3a",  x"41",  x"03",  x"47", -- 06E0
         x"3a",  x"ac",  x"31",  x"03",  x"04",  x"ba",  x"06",  x"05", -- 06E8
         x"b8",  x"cc",  x"61",  x"cb",  x"88",  x"5a",  x"0b",  x"79", -- 06F0
         x"80",  x"d4",  x"c1",  x"f1",  x"6b",  x"c9",  x"e7",  x"a6", -- 06F8
         x"b7",  x"2e",  x"09",  x"af",  x"04",  x"7b",  x"3c",  x"69", -- 0700
         x"4a",  x"fd",  x"b1",  x"d3",  x"22",  x"61",  x"8c",  x"64", -- 0708
         x"63",  x"03",  x"65",  x"82",  x"41",  x"6c",  x"c9",  x"ed", -- 0710
         x"53",  x"46",  x"da",  x"68",  x"89",  x"80",  x"25",  x"de", -- 0718
         x"cd",  x"c8",  x"dd",  x"28",  x"12",  x"90",  x"c5",  x"1d", -- 0720
         x"2a",  x"13",  x"ab",  x"a6",  x"ff",  x"b4",  x"cd",  x"08", -- 0728
         x"e1",  x"3a",  x"a3",  x"80",  x"c5",  x"cd",  x"91",  x"c7", -- 0730
         x"e1",  x"4e",  x"23",  x"00",  x"46",  x"23",  x"78",  x"b1", -- 0738
         x"28",  x"59",  x"cd",  x"67",  x"00",  x"c7",  x"cd",  x"f9", -- 0740
         x"c8",  x"c5",  x"5e",  x"23",  x"56",  x"29",  x"23",  x"e5", -- 0748
         x"8f",  x"9d",  x"cd",  x"71",  x"36",  x"84",  x"8f",  x"1f", -- 0750
         x"2c",  x"65",  x"9e",  x"ee",  x"d2",  x"66",  x"28",  x"14", -- 0758
         x"b9",  x"43",  x"d3",  x"f2",  x"3c",  x"23",  x"7b",  x"9a", -- 0760
         x"02",  x"11",  x"1a",  x"cb",  x"40",  x"f2",  x"4e",  x"c7", -- 0768
         x"18",  x"49",  x"e6",  x"1c",  x"a8",  x"18",  x"ba",  x"1f", -- 0770
         x"d7",  x"18",  x"6e",  x"f2",  x"bf",  x"44",  x"63",  x"03", -- 0778
         x"d2",  x"8e",  x"9a",  x"05",  x"e1",  x"55",  x"c0",  x"5a", -- 0780
         x"10",  x"c2",  x"fe",  x"03",  x"20",  x"58",  x"ea",  x"84", -- 0788
         x"2f",  x"0c",  x"4e",  x"ee",  x"66",  x"2a",  x"82",  x"15", -- 0790
         x"7f",  x"5d",  x"8b",  x"f6",  x"29",  x"06",  x"26",  x"c9", -- 0798
         x"0d",  x"d6",  x"7f",  x"fe",  x"56",  x"d7",  x"4c",  x"d6", -- 07A0
         x"55",  x"96",  x"b3",  x"e3",  x"6e",  x"18",  x"b0",  x"21", -- 07A8
         x"2c",  x"c1",  x"47",  x"5a",  x"ac",  x"c7",  x"33",  x"10", -- 07B0
         x"f8",  x"f0",  x"56",  x"c9",  x"be",  x"b0",  x"0a",  x"ca", -- 07B8
         x"78",  x"21",  x"a0",  x"39",  x"a0",  x"81",  x"2c",  x"81", -- 07C0
         x"c0",  x"a9",  x"00",  x"e5",  x"69",  x"60",  x"7a",  x"b3", -- 07C8
         x"eb",  x"cd",  x"d8",  x"eb",  x"42",  x"b0",  x"01",  x"e0", -- 07D0
         x"b7",  x"e1",  x"c8",  x"05",  x"09",  x"18",  x"e3",  x"3e", -- 07D8
         x"64",  x"0b",  x"e2",  x"cd",  x"95",  x"a6",  x"c1",  x"f8", -- 07E0
         x"bd",  x"a2",  x"18",  x"22",  x"c8",  x"e5",  x"30",  x"02", -- 07E8
         x"30",  x"cd",  x"c1",  x"c7",  x"d1",  x"cc",  x"ab",  x"09", -- 07F0
         x"d5",  x"18",  x"2b",  x"56",  x"2b",  x"d1",  x"6e",  x"35", -- 07F8
         x"2a",  x"15",  x"80",  x"30",  x"e1",  x"20",  x"e8",  x"d1", -- 0800
         x"f9",  x"eb",  x"33",  x"0e",  x"08",  x"a7",  x"5b",  x"c3", -- 0808
         x"11",  x"e3",  x"04",  x"7f",  x"58",  x"04",  x"b4",  x"00", -- 0810
         x"cd",  x"cd",  x"cc",  x"c8",  x"a6",  x"cd",  x"26",  x"60", -- 0818
         x"cd",  x"3e",  x"eb",  x"d6",  x"e1",  x"c5",  x"d5",  x"06", -- 0820
         x"01",  x"00",  x"81",  x"51",  x"5a",  x"a2",  x"40",  x"ab", -- 0828
         x"3e",  x"01",  x"20",  x"0e",  x"a4",  x"e1",  x"9b",  x"18", -- 0830
         x"d0",  x"1b",  x"1b",  x"36",  x"f5",  x"33",  x"33",  x"cf", -- 0838
         x"33",  x"06",  x"02",  x"81",  x"c5",  x"33",  x"cd",  x"16", -- 0840
         x"de",  x"86",  x"af",  x"8f",  x"86",  x"2a",  x"d0",  x"e8", -- 0848
         x"28",  x"b7",  x"a3",  x"ce",  x"a6",  x"9f",  x"65",  x"b6", -- 0850
         x"7f",  x"c9",  x"23",  x"0e",  x"c2",  x"83",  x"59",  x"59", -- 0858
         x"3a",  x"0a",  x"50",  x"d1",  x"0f",  x"e5",  x"ca",  x"3c", -- 0860
         x"65",  x"a7",  x"43",  x"ca",  x"6e",  x"ef",  x"e1",  x"a3", -- 0868
         x"50",  x"11",  x"54",  x"d7",  x"70",  x"c8",  x"d6",  x"80", -- 0870
         x"da",  x"c0",  x"b0",  x"fe",  x"25",  x"00",  x"38",  x"14", -- 0878
         x"d6",  x"50",  x"38",  x"34",  x"fe",  x"05",  x"16",  x"38", -- 0880
         x"0a",  x"47",  x"f2",  x"a0",  x"28",  x"29",  x"c3",  x"03", -- 0888
         x"e0",  x"0e",  x"c6",  x"25",  x"07",  x"4f",  x"85",  x"b7", -- 0890
         x"a4",  x"14",  x"40",  x"c2",  x"09",  x"f1",  x"0d",  x"c5", -- 0898
         x"96",  x"a9",  x"60",  x"d0",  x"99",  x"90",  x"28",  x"f7", -- 08A0
         x"b3",  x"c0",  x"3f",  x"a3",  x"8c",  x"bc",  x"db",  x"e3", -- 08A8
         x"ac",  x"e8",  x"cb",  x"ea",  x"63",  x"c3",  x"6f",  x"3e", -- 08B0
         x"2c",  x"be",  x"9f",  x"71",  x"3e",  x"29",  x"18",  x"85", -- 08B8
         x"d2",  x"26",  x"90",  x"a6",  x"aa",  x"eb",  x"d6",  x"25", -- 08C0
         x"e5",  x"16",  x"d5",  x"9e",  x"e6",  x"d1",  x"d2",  x"87", -- 08C8
         x"f9",  x"85",  x"38",  x"dd",  x"80",  x"cc",  x"86",  x"f3", -- 08D0
         x"dd",  x"06",  x"c0",  x"fe",  x"13",  x"28",  x"08",  x"87", -- 08D8
         x"4a",  x"c0",  x"8d",  x"22",  x"18",  x"0f",  x"c8",  x"92", -- 08E0
         x"1e",  x"c8",  x"3c",  x"fe",  x"0a",  x"02",  x"30",  x"02", -- 08E8
         x"18",  x"0a",  x"f1",  x"c0",  x"f6",  x"c0",  x"c0",  x"00", -- 08F0
         x"21",  x"f6",  x"ff",  x"c1",  x"a1",  x"89",  x"0d",  x"f5", -- 08F8
         x"7d",  x"a4",  x"3c",  x"9c",  x"8d",  x"22",  x"d3",  x"d7", -- 0900
         x"3a",  x"12",  x"b6",  x"49",  x"2b",  x"ab",  x"c3",  x"4a", -- 0908
         x"ae",  x"a0",  x"f1",  x"21",  x"21",  x"c3",  x"01",  x"c2", -- 0910
         x"71",  x"c3",  x"c3",  x"88",  x"c3",  x"2a",  x"8c",  x"16", -- 0918
         x"7c",  x"b5",  x"1e",  x"5c",  x"56",  x"c3",  x"d7",  x"72", -- 0920
         x"d3",  x"90",  x"7c",  x"61",  x"a3",  x"a1",  x"42",  x"9d", -- 0928
         x"f2",  x"07",  x"6f",  x"c9",  x"1e",  x"08",  x"c3",  x"19", -- 0930
         x"40",  x"0d",  x"3a",  x"e8",  x"03",  x"fe",  x"90",  x"01", -- 0938
         x"da",  x"45",  x"d7",  x"01",  x"80",  x"90",  x"11",  x"fe", -- 0940
         x"db",  x"93",  x"00",  x"18",  x"d7",  x"e1",  x"51",  x"c8", -- 0948
         x"15",  x"18",  x"e1",  x"2b",  x"0c",  x"40",  x"2e",  x"d0", -- 0950
         x"e5",  x"f5",  x"21",  x"98",  x"51",  x"19",  x"8e",  x"30", -- 0958
         x"da",  x"c2",  x"e4",  x"85",  x"19",  x"29",  x"c0",  x"01", -- 0960
         x"f1",  x"d6",  x"30",  x"5f",  x"16",  x"00",  x"37",  x"19", -- 0968
         x"eb",  x"c0",  x"31",  x"e0",  x"28",  x"ad",  x"62",  x"5e", -- 0970
         x"53",  x"be",  x"c8",  x"e5",  x"94",  x"dc",  x"28",  x"10", -- 0978
         x"53",  x"e1",  x"b0",  x"68",  x"bd",  x"6c",  x"ba",  x"10", -- 0980
         x"df",  x"16",  x"e3",  x"af",  x"c0",  x"93",  x"5f",  x"7c", -- 0988
         x"9a",  x"57",  x"28",  x"da",  x"3e",  x"be",  x"b5",  x"f1", -- 0990
         x"3c",  x"01",  x"28",  x"aa",  x"a6",  x"45",  x"d2",  x"0d", -- 0998
         x"eb",  x"29",  x"22",  x"56",  x"bd",  x"bd",  x"30",  x"8a", -- 09A0
         x"dd",  x"53",  x"ed",  x"f2",  x"e0",  x"cd",  x"cc",  x"05", -- 09A8
         x"01",  x"54",  x"6f",  x"10",  x"0e",  x"51",  x"03",  x"e8", -- 09B0
         x"67",  x"94",  x"21",  x"e5",  x"19",  x"3e",  x"8c",  x"ba", -- 09B8
         x"68",  x"ee",  x"86",  x"fd",  x"49",  x"f8",  x"bb",  x"0f", -- 09C0
         x"8c",  x"30",  x"23",  x"dc",  x"be",  x"c4",  x"58",  x"d4", -- 09C8
         x"ae",  x"bc",  x"2b",  x"e1",  x"50",  x"0e",  x"b8",  x"1d", -- 09D0
         x"c0",  x"16",  x"cf",  x"80",  x"bd",  x"c7",  x"f9",  x"fe", -- 09D8
         x"8c",  x"1e",  x"04",  x"3d",  x"20",  x"f0",  x"4e",  x"24", -- 09E0
         x"23",  x"80",  x"eb",  x"20",  x"07",  x"3a",  x"eb",  x"ff", -- 09E8
         x"db",  x"27",  x"87",  x"a2",  x"7e",  x"50",  x"43",  x"e1", -- 09F0
         x"0c",  x"01",  x"3a",  x"0e",  x"00",  x"9a",  x"8a",  x"79", -- 09F8
         x"48",  x"c6",  x"81",  x"c8",  x"b8",  x"c8",  x"6a",  x"95", -- 0A00
         x"f3",  x"05",  x"18",  x"f4",  x"cd",  x"06",  x"cf",  x"18", -- 0A08
         x"c0",  x"b4",  x"d5",  x"3a",  x"62",  x"ae",  x"c2",  x"cd", -- 0A10
         x"ca",  x"2e",  x"f1",  x"e3",  x"d2",  x"10",  x"1f",  x"cd", -- 0A18
         x"2b",  x"cd",  x"36",  x"28",  x"35",  x"69",  x"e5",  x"f7", -- 0A20
         x"cb",  x"23",  x"8f",  x"3c",  x"a0",  x"ac",  x"72",  x"30", -- 0A28
         x"12",  x"a7",  x"9e",  x"93",  x"b3",  x"34",  x"e8",  x"49", -- 0A30
         x"c0",  x"10",  x"e8",  x"ea",  x"d1",  x"cd",  x"1b",  x"64", -- 0A38
         x"d3",  x"b9",  x"66",  x"bc",  x"06",  x"ed",  x"19",  x"fa", -- 0A40
         x"e3",  x"d1",  x"c2",  x"3d",  x"f7",  x"c2",  x"a8",  x"cb", -- 0A48
         x"1d",  x"21",  x"d4",  x"7e",  x"c9",  x"36",  x"8c",  x"fc", -- 0A50
         x"a3",  x"5b",  x"88",  x"2b",  x"a2",  x"e1",  x"78",  x"ca", -- 0A58
         x"92",  x"88",  x"e8",  x"87",  x"c9",  x"fe",  x"39",  x"2c", -- 0A60
         x"c0",  x"b7",  x"ac",  x"65",  x"93",  x"d2",  x"88",  x"35", -- 0A68
         x"1a",  x"a9",  x"67",  x"29",  x"88",  x"fd",  x"20",  x"08", -- 0A70
         x"23",  x"a0",  x"93",  x"0a",  x"fe",  x"d4",  x"20",  x"f8", -- 0A78
         x"e1",  x"10",  x"da",  x"07",  x"ca",  x"c3",  x"78",  x"91", -- 0A80
         x"2d",  x"b4",  x"99",  x"18",  x"07",  x"c5",  x"3d",  x"fd", -- 0A88
         x"68",  x"88",  x"cc",  x"28",  x"5e",  x"1b",  x"d5",  x"38", -- 0A90
         x"48",  x"09",  x"e3",  x"78",  x"0f",  x"06",  x"e0",  x"fe", -- 0A98
         x"60",  x"a5",  x"4e",  x"cb",  x"fe",  x"a8",  x"28",  x"78", -- 0AA0
         x"60",  x"e5",  x"50",  x"28",  x"5d",  x"fe",  x"3b",  x"ca", -- 0AA8
         x"14",  x"b2",  x"cb",  x"c1",  x"55",  x"e5",  x"a0",  x"c3", -- 0AB0
         x"f3",  x"a4",  x"ef",  x"d0",  x"34",  x"d8",  x"cd",  x"8a", -- 0AB8
         x"14",  x"d1",  x"36",  x"20",  x"be",  x"0a",  x"34",  x"03", -- 0AC0
         x"b8",  x"88",  x"e0",  x"85",  x"0a",  x"04",  x"a8",  x"8c", -- 0AC8
         x"0d",  x"86",  x"3d",  x"b8",  x"d4",  x"c9",  x"bc",  x"77", -- 0AD0
         x"a0",  x"0f",  x"18",  x"a0",  x"0e",  x"2b",  x"c5",  x"61", -- 0AD8
         x"05",  x"36",  x"00",  x"51",  x"91",  x"3e",  x"0d",  x"70", -- 0AE0
         x"91",  x"0a",  x"af",  x"04",  x"70",  x"16",  x"01",  x"3a", -- 0AE8
         x"40",  x"03",  x"3d",  x"c8",  x"f5",  x"af",  x"4d",  x"0d", -- 0AF0
         x"f1",  x"a0",  x"09",  x"3a",  x"42",  x"22",  x"c6",  x"c3", -- 0AF8
         x"37",  x"30",  x"29",  x"d6",  x"0d",  x"ab",  x"b0",  x"20", -- 0B00
         x"fa",  x"2f",  x"18",  x"62",  x"15",  x"a9",  x"1e",  x"1d", -- 0B08
         x"d4",  x"cd",  x"db",  x"be",  x"e4",  x"fa",  x"a8",  x"61", -- 0B10
         x"e5",  x"91",  x"41",  x"1f",  x"2f",  x"83",  x"30",  x"0b", -- 0B18
         x"99",  x"fe",  x"08",  x"47",  x"27",  x"ed",  x"16",  x"10", -- 0B20
         x"fb",  x"a8",  x"ba",  x"8b",  x"f8",  x"69",  x"85",  x"bb", -- 0B28
         x"32",  x"7d",  x"8c",  x"1a",  x"88",  x"cc",  x"55",  x"c9", -- 0B30
         x"3f",  x"00",  x"52",  x"45",  x"44",  x"4f",  x"20",  x"46", -- 0B38
         x"52",  x"4f",  x"3b",  x"4d",  x"20",  x"b1",  x"1b",  x"41", -- 0B40
         x"52",  x"54",  x"81",  x"94",  x"3a",  x"ce",  x"9f",  x"4c", -- 0B48
         x"42",  x"e6",  x"8f",  x"21",  x"c9",  x"2c",  x"d3",  x"f3", -- 0B50
         x"c3",  x"85",  x"fd",  x"22",  x"37",  x"d1",  x"aa",  x"c1", -- 0B58
         x"d3",  x"bd",  x"a3",  x"10",  x"22",  x"20",  x"10",  x"cd", -- 0B60
         x"78",  x"8b",  x"0e",  x"a6",  x"9e",  x"3b",  x"e5",  x"04", -- 0B68
         x"07",  x"d4",  x"18",  x"c6",  x"18",  x"04",  x"08",  x"cf", -- 0B70
         x"c6",  x"c1",  x"2a",  x"38",  x"36",  x"bb",  x"f1",  x"af", -- 0B78
         x"76",  x"2b",  x"d5",  x"37",  x"30",  x"36",  x"2c",  x"c2", -- 0B80
         x"cb",  x"a7",  x"ab",  x"57",  x"f6",  x"31",  x"b8",  x"49", -- 0B88
         x"e3",  x"82",  x"a3",  x"f1",  x"a2",  x"d0",  x"7f",  x"e3", -- 0B90
         x"bc",  x"42",  x"98",  x"1e",  x"b2",  x"5c",  x"20",  x"7d", -- 0B98
         x"49",  x"ee",  x"a0",  x"36",  x"d1",  x"c1",  x"da",  x"1f", -- 0BA0
         x"4c",  x"c9",  x"38",  x"ca",  x"2c",  x"47",  x"ca",  x"f0", -- 0BA8
         x"b6",  x"e0",  x"50",  x"21",  x"a8",  x"2b",  x"57",  x"f2", -- 0BB0
         x"78",  x"e2",  x"b6",  x"2c",  x"57",  x"d5",  x"a1",  x"16", -- 0BB8
         x"3a",  x"06",  x"2c",  x"91",  x"94",  x"8e",  x"d1",  x"b1", -- 0BC0
         x"c0",  x"88",  x"cc",  x"8b",  x"46",  x"c3",  x"77",  x"ca", -- 0BC8
         x"a1",  x"51",  x"a1",  x"d7",  x"e3",  x"44",  x"d6",  x"e1", -- 0BD0
         x"a2",  x"92",  x"cb",  x"b5",  x"58",  x"1e",  x"c2",  x"db", -- 0BD8
         x"cb",  x"0e",  x"0a",  x"20",  x"2c",  x"93",  x"d1",  x"33", -- 0BE0
         x"eb",  x"c2",  x"68",  x"f4",  x"e4",  x"b6",  x"05",  x"21", -- 0BE8
         x"ab",  x"cc",  x"c4",  x"c9",  x"10",  x"f7",  x"3f",  x"45", -- 0BF0
         x"58",  x"00",  x"54",  x"52",  x"41",  x"20",  x"49",  x"47", -- 0BF8
         x"4e",  x"4f",  x"a0",  x"eb",  x"c2",  x"df",  x"a3",  x"d2", -- 0C00
         x"82",  x"05",  x"11",  x"b9",  x"da",  x"1e",  x"06",  x"4b", -- 0C08
         x"f7",  x"2b",  x"dc",  x"94",  x"ca",  x"03",  x"54",  x"fe", -- 0C10
         x"1a",  x"83",  x"20",  x"e2",  x"b6",  x"29",  x"cc",  x"d4", -- 0C18
         x"58",  x"c4",  x"b0",  x"51",  x"f3",  x"d2",  x"bc",  x"03", -- 0C20
         x"c2",  x"4e",  x"c3",  x"f9",  x"d5",  x"2a",  x"6a",  x"f5", -- 0C28
         x"b3",  x"dd",  x"71",  x"d6",  x"dd",  x"cb",  x"f3",  x"d4", -- 0C30
         x"71",  x"b2",  x"75",  x"ee",  x"d6",  x"46",  x"83",  x"2b", -- 0C38
         x"c1",  x"90",  x"09",  x"e1",  x"6b",  x"9b",  x"8e",  x"c5", -- 0C40
         x"41",  x"c3",  x"50",  x"c8",  x"f9",  x"2a",  x"71",  x"bc", -- 0C48
         x"86",  x"8d",  x"da",  x"96",  x"a2",  x"05",  x"df",  x"cc", -- 0C50
         x"19",  x"80",  x"f6",  x"37",  x"40",  x"d4",  x"8f",  x"0b", -- 0C58
         x"b7",  x"e8",  x"1e",  x"18",  x"c9",  x"6c",  x"b7",  x"4d", -- 0C60
         x"28",  x"2b",  x"97",  x"86",  x"d5",  x"0e",  x"01",  x"c7", -- 0C68
         x"b8",  x"0c",  x"ad",  x"cd",  x"22",  x"6f",  x"d1",  x"9a", -- 0C70
         x"be",  x"02",  x"c1",  x"fa",  x"33",  x"78",  x"d4",  x"f3", -- 0C78
         x"61",  x"7e",  x"18",  x"d6",  x"b3",  x"38",  x"15",  x"be", -- 0C80
         x"c7",  x"cb",  x"80",  x"fe",  x"01",  x"17",  x"aa",  x"ba", -- 0C88
         x"53",  x"57",  x"cd",  x"16",  x"22",  x"c6",  x"97",  x"03", -- 0C90
         x"18",  x"e7",  x"7a",  x"91",  x"21",  x"84",  x"ce",  x"7e", -- 0C98
         x"47",  x"0d",  x"d6",  x"ac",  x"e7",  x"82",  x"07",  x"d0", -- 0CA0
         x"5f",  x"80",  x"53",  x"3d",  x"b3",  x"7b",  x"ca",  x"b3", -- 0CA8
         x"d2",  x"0d",  x"07",  x"83",  x"5f",  x"21",  x"c9",  x"80", -- 0CB0
         x"19",  x"78",  x"56",  x"ba",  x"d0",  x"23",  x"a4",  x"b7", -- 0CB8
         x"19",  x"c5",  x"01",  x"49",  x"03",  x"43",  x"4a",  x"d8", -- 0CC0
         x"a0",  x"d6",  x"58",  x"51",  x"ba",  x"dc",  x"f7",  x"a2", -- 0CC8
         x"32",  x"32",  x"18",  x"90",  x"88",  x"59",  x"ae",  x"46", -- 0CD0
         x"1e",  x"24",  x"40",  x"ee",  x"da",  x"c4",  x"b8",  x"cd", -- 0CD8
         x"8f",  x"d4",  x"a6",  x"37",  x"fe",  x"03",  x"ac",  x"28", -- 0CE0
         x"e8",  x"fe",  x"2e",  x"ca",  x"0d",  x"0c",  x"fe",  x"ad", -- 0CE8
         x"28",  x"19",  x"ec",  x"59",  x"ca",  x"d4",  x"00",  x"fe", -- 0CF0
         x"aa",  x"ca",  x"e3",  x"ce",  x"fe",  x"a7",  x"00",  x"ca", -- 0CF8
         x"f0",  x"d0",  x"d6",  x"b6",  x"30",  x"28",  x"cd",  x"19", -- 0D00
         x"36",  x"cd",  x"c3",  x"cd",  x"82",  x"16",  x"7d",  x"cd", -- 0D08
         x"3d",  x"cd",  x"83",  x"a2",  x"ed",  x"02",  x"c0",  x"d6", -- 0D10
         x"a9",  x"5e",  x"c4",  x"71",  x"98",  x"6f",  x"e5",  x"9c", -- 0D18
         x"a5",  x"c1",  x"93",  x"a9",  x"cc",  x"92",  x"1f",  x"10", -- 0D20
         x"bc",  x"6e",  x"db",  x"54",  x"c5",  x"5c",  x"79",  x"0b", -- 0D28
         x"fe",  x"33",  x"38",  x"07",  x"8d",  x"5e",  x"e3",  x"5e", -- 0D30
         x"e0",  x"4e",  x"e8",  x"41",  x"fe",  x"2d",  x"38",  x"17", -- 0D38
         x"56",  x"43",  x"fc",  x"4e",  x"2a",  x"ec",  x"a9",  x"f3", -- 0D40
         x"1d",  x"e3",  x"37",  x"1f",  x"f4",  x"b4",  x"e6",  x"18", -- 0D48
         x"08",  x"46",  x"cd",  x"35",  x"e3",  x"11",  x"f2",  x"ed", -- 0D50
         x"96",  x"94",  x"74",  x"8f",  x"66",  x"30",  x"69",  x"e9", -- 0D58
         x"f3",  x"30",  x"ad",  x"c8",  x"2f",  x"c8",  x"14",  x"fe", -- 0D60
         x"2b",  x"da",  x"06",  x"ac",  x"c1",  x"33",  x"c9",  x"b9", -- 0D68
         x"5b",  x"f5",  x"83",  x"70",  x"fe",  x"f1",  x"18",  x"eb", -- 0D70
         x"c1",  x"e3",  x"35",  x"e0",  x"d6",  x"f5",  x"b0",  x"0b", -- 0D78
         x"c1",  x"79",  x"21",  x"b0",  x"00",  x"d0",  x"20",  x"05", -- 0D80
         x"a3",  x"4f",  x"78",  x"a2",  x"e9",  x"60",  x"b3",  x"04", -- 0D88
         x"b2",  x"e9",  x"21",  x"96",  x"ce",  x"a0",  x"86",  x"1c", -- 0D90
         x"1f",  x"7a",  x"17",  x"ea",  x"18",  x"64",  x"78",  x"ff", -- 0D98
         x"00",  x"c3",  x"97",  x"cd",  x"98",  x"ce",  x"79",  x"b7", -- 0DA0
         x"1b",  x"1f",  x"c1",  x"d1",  x"2e",  x"2b",  x"6a",  x"0c", -- 0DA8
         x"d9",  x"ce",  x"e5",  x"ca",  x"a2",  x"ac",  x"fa",  x"32", -- 0DB0
         x"bb",  x"32",  x"fe",  x"d2",  x"c2",  x"50",  x"23",  x"8f", -- 0DB8
         x"99",  x"d1",  x"c5",  x"1a",  x"02",  x"d3",  x"44",  x"b3", -- 0DC0
         x"f1",  x"00",  x"57",  x"e1",  x"7b",  x"b2",  x"c8",  x"7a", -- 0DC8
         x"d6",  x"01",  x"00",  x"d8",  x"af",  x"bb",  x"3c",  x"d0", -- 0DD0
         x"15",  x"1d",  x"0a",  x"ef",  x"81",  x"9c",  x"90",  x"ed", -- 0DD8
         x"3f",  x"c3",  x"a2",  x"00",  x"d6",  x"3c",  x"8f",  x"c1", -- 0DE0
         x"a0",  x"c6",  x"ff",  x"9f",  x"05",  x"c3",  x"a9",  x"d6", -- 0DE8
         x"16",  x"5a",  x"04",  x"fb",  x"a0",  x"87",  x"7b",  x"06", -- 0DF0
         x"2f",  x"4f",  x"7a",  x"2f",  x"cd",  x"7d",  x"c1",  x"63", -- 0DF8
         x"c3",  x"de",  x"46",  x"e6",  x"c8",  x"a0",  x"d5",  x"0a", -- 0E00
         x"01",  x"fa",  x"ce",  x"c5",  x"e1",  x"41",  x"ad",  x"03", -- 0E08
         x"46",  x"8d",  x"ce",  x"c9",  x"f7",  x"af",  x"4f",  x"28", -- 0E10
         x"e4",  x"94",  x"38",  x"05",  x"0f",  x"38",  x"2d",  x"0b", -- 0E18
         x"4f",  x"0a",  x"fb",  x"62",  x"e9",  x"f6",  x"05",  x"d6", -- 0E20
         x"24",  x"20",  x"0a",  x"3c",  x"16",  x"1c",  x"0f",  x"81", -- 0E28
         x"14",  x"3a",  x"f4",  x"d8",  x"3d",  x"ca",  x"03",  x"dd", -- 0E30
         x"cf",  x"f2",  x"48",  x"cf",  x"7e",  x"b9",  x"33",  x"28", -- 0E38
         x"6f",  x"41",  x"c1",  x"0f",  x"e5",  x"50",  x"59",  x"2a", -- 0E40
         x"df",  x"70",  x"bc",  x"11",  x"01",  x"e1",  x"03",  x"ca", -- 0E48
         x"e0",  x"d5",  x"2a",  x"d9",  x"df",  x"84",  x"8c",  x"57", -- 0E50
         x"0f",  x"d0",  x"ae",  x"79",  x"96",  x"23",  x"18",  x"20", -- 0E58
         x"02",  x"78",  x"04",  x"28",  x"38",  x"23",  x"a7",  x"00", -- 0E60
         x"18",  x"cf",  x"5a",  x"ff",  x"3b",  x"11",  x"55",  x"f0", -- 0E68
         x"8f",  x"d8",  x"31",  x"d0",  x"cb",  x"ed",  x"fd",  x"13", -- 0E70
         x"2a",  x"db",  x"3f",  x"57",  x"09",  x"a7",  x"1c",  x"ab", -- 0E78
         x"c4",  x"e0",  x"fc",  x"0a",  x"fa",  x"b6",  x"22",  x"3d", -- 0E80
         x"2b",  x"c0",  x"f5",  x"21",  x"c0",  x"b7",  x"d1",  x"73", -- 0E88
         x"23",  x"33",  x"72",  x"23",  x"32",  x"c9",  x"32",  x"bc", -- 0E90
         x"b1",  x"21",  x"20",  x"c3",  x"45",  x"b4",  x"ed",  x"0a", -- 0E98
         x"97",  x"80",  x"b0",  x"e3",  x"57",  x"d5",  x"c8",  x"b0", -- 0EA0
         x"5b",  x"c9",  x"63",  x"c1",  x"dc",  x"44",  x"92",  x"3c", -- 0EA8
         x"5b",  x"57",  x"96",  x"29",  x"ee",  x"b8",  x"e9",  x"8b", -- 0EB0
         x"3c",  x"41",  x"1d",  x"1e",  x"00",  x"fb",  x"61",  x"ce", -- 0EB8
         x"a0",  x"83",  x"3f",  x"3e",  x"19",  x"c1",  x"ec",  x"50", -- 0EC0
         x"85",  x"35",  x"aa",  x"50",  x"b9",  x"85",  x"16",  x"7e", -- 0EC8
         x"b8",  x"a9",  x"b9",  x"08",  x"e8",  x"3a",  x"e8",  x"24", -- 0ED0
         x"8d",  x"51",  x"00",  x"c3",  x"f1",  x"44",  x"4d",  x"ca", -- 0ED8
         x"aa",  x"cf",  x"96",  x"0a",  x"28",  x"5f",  x"1e",  x"10", -- 0EE0
         x"d9",  x"47",  x"11",  x"d2",  x"e0",  x"f1",  x"ca",  x"67", -- 0EE8
         x"c9",  x"71",  x"0a",  x"23",  x"70",  x"23",  x"4f",  x"db", -- 0EF0
         x"4c",  x"ab",  x"29",  x"ab",  x"3a",  x"0c",  x"2a",  x"00", -- 0EF8
         x"17",  x"79",  x"01",  x"0b",  x"00",  x"30",  x"02",  x"c1", -- 0F00
         x"59",  x"03",  x"1a",  x"f5",  x"e5",  x"b0",  x"4f",  x"d7", -- 0F08
         x"91",  x"00",  x"f1",  x"3d",  x"20",  x"ea",  x"f5",  x"42", -- 0F10
         x"4b",  x"eb",  x"55",  x"19",  x"f7",  x"98",  x"cd",  x"30", -- 0F18
         x"99",  x"73",  x"66",  x"81",  x"b2",  x"03",  x"57",  x"48", -- 0F20
         x"b0",  x"5e",  x"02",  x"eb",  x"29",  x"09",  x"eb",  x"2b", -- 0F28
         x"2b",  x"c0",  x"bd",  x"f1",  x"38",  x"19",  x"22",  x"47", -- 0F30
         x"4f",  x"bb",  x"16",  x"16",  x"e1",  x"7a",  x"e3",  x"5d", -- 0F38
         x"f5",  x"e0",  x"2c",  x"90",  x"43",  x"d1",  x"19",  x"fc", -- 0F40
         x"43",  x"7f",  x"8b",  x"07",  x"29",  x"29",  x"c1",  x"2a", -- 0F48
         x"48",  x"9f",  x"c9",  x"b0",  x"ab",  x"6c",  x"21",  x"b7", -- 0F50
         x"39",  x"91",  x"c1",  x"d4",  x"0d",  x"f0",  x"43",  x"cd", -- 0F58
         x"09",  x"d2",  x"13",  x"ec",  x"9b",  x"2a",  x"c4",  x"78", -- 0F60
         x"03",  x"e2",  x"4f",  x"f0",  x"e2",  x"41",  x"50",  x"c1", -- 0F68
         x"d8",  x"21",  x"81",  x"1b",  x"73",  x"06",  x"90",  x"c3", -- 0F70
         x"ae",  x"d6",  x"52",  x"9c",  x"47",  x"02",  x"af",  x"18", -- 0F78
         x"ed",  x"cd",  x"45",  x"d1",  x"a1",  x"da",  x"01",  x"b9", -- 0F80
         x"8e",  x"c5",  x"d5",  x"6d",  x"98",  x"69",  x"da",  x"85", -- 0F88
         x"76",  x"56",  x"2b",  x"5e",  x"e1",  x"96",  x"f4",  x"90", -- 0F90
         x"37",  x"82",  x"9a",  x"63",  x"e3",  x"80",  x"b7",  x"c3", -- 0F98
         x"84",  x"ff",  x"28",  x"2b",  x"24",  x"18",  x"a5",  x"19", -- 0FA0
         x"e3",  x"80",  x"8a",  x"7a",  x"b3",  x"ca",  x"30",  x"54", -- 0FA8
         x"c3",  x"97",  x"14",  x"66",  x"6f",  x"e5",  x"b9",  x"5e", -- 0FB0
         x"9e",  x"63",  x"03",  x"2a",  x"e3",  x"03",  x"0a",  x"6f", -- 0FB8
         x"e1",  x"03",  x"21",  x"03",  x"27",  x"b7",  x"a1",  x"fa", -- 0FC0
         x"b3",  x"5d",  x"e2",  x"c7",  x"d3",  x"11",  x"ff",  x"03", -- 0FC8
         x"1d",  x"03",  x"24",  x"b1",  x"ff",  x"93",  x"84",  x"42", -- 0FD0
         x"e1",  x"c0",  x"1e",  x"16",  x"57",  x"8e",  x"14",  x"a7", -- 0FD8
         x"3e",  x"80",  x"81",  x"60",  x"b6",  x"47",  x"cd",  x"0b", -- 0FE0
         x"cf",  x"2e",  x"c3",  x"29",  x"5e",  x"5b",  x"a9",  x"a0", -- 0FE8
         x"c0",  x"0a",  x"01",  x"57",  x"d3",  x"c5",  x"b5",  x"47", -- 0FF0
         x"e5",  x"75",  x"c5",  x"c3",  x"26",  x"ba",  x"9e",  x"e0", -- 0FF8
         x"d1",  x"e5",  x"6f",  x"cd",  x"f2",  x"15",  x"d2",  x"d1", -- 1000
         x"c9",  x"10",  x"e6",  x"eb",  x"69",  x"77",  x"e8",  x"1b", -- 1008
         x"a1",  x"70",  x"52",  x"2b",  x"06",  x"22",  x"50",  x"19", -- 1010
         x"e5",  x"0e",  x"ff",  x"a4",  x"30",  x"0c",  x"f8",  x"3a", -- 1018
         x"06",  x"ba",  x"f9",  x"1a",  x"b8",  x"20",  x"f4",  x"ff", -- 1020
         x"b3",  x"cc",  x"e8",  x"64",  x"e3",  x"fa",  x"79",  x"a6", -- 1028
         x"34",  x"11",  x"2a",  x"2a",  x"28",  x"b2",  x"03",  x"fc", -- 1030
         x"8b",  x"3e",  x"01",  x"a0",  x"4f",  x"8f",  x"68",  x"c3", -- 1038
         x"59",  x"22",  x"10",  x"e1",  x"7e",  x"82",  x"82",  x"1e", -- 1040
         x"81",  x"82",  x"23",  x"2d",  x"6c",  x"28",  x"92",  x"1c", -- 1048
         x"1d",  x"c8",  x"bb",  x"ed",  x"06",  x"fe",  x"0d",  x"cc", -- 1050
         x"66",  x"cb",  x"b3",  x"e0",  x"f2",  x"b7",  x"0e",  x"f1", -- 1058
         x"f5",  x"98",  x"c0",  x"74",  x"fc",  x"1f",  x"06",  x"ff", -- 1060
         x"09",  x"28",  x"37",  x"b3",  x"e0",  x"22",  x"0d",  x"db", -- 1068
         x"56",  x"f1",  x"8b",  x"00",  x"1e",  x"1a",  x"28",  x"c2", -- 1070
         x"bf",  x"f5",  x"01",  x"6b",  x"e3",  x"d0",  x"5f",  x"d5", -- 1078
         x"d8",  x"14",  x"fa",  x"e1",  x"da",  x"e0",  x"2c",  x"fe", -- 1080
         x"b4",  x"7d",  x"03",  x"34",  x"5d",  x"02",  x"2b",  x"01", -- 1088
         x"1a",  x"d2",  x"20",  x"3f",  x"93",  x"c6",  x"0e",  x"5f", -- 1090
         x"d9",  x"0e",  x"ec",  x"94",  x"cb",  x"00",  x"b7",  x"cd", -- 1098
         x"68",  x"d2",  x"18",  x"27",  x"ee",  x"c1",  x"d7",  x"35", -- 10A0
         x"49",  x"34",  x"75",  x"7b",  x"bc",  x"0a",  x"b7",  x"f2", -- 10A8
         x"3b",  x"d2",  x"ad",  x"3c",  x"e4",  x"34",  x"cc",  x"7f", -- 10B0
         x"09",  x"66",  x"1c",  x"0a",  x"61",  x"1c",  x"da",  x"01", -- 10B8
         x"59",  x"d2",  x"aa",  x"e0",  x"80",  x"ac",  x"35",  x"ef", -- 10C0
         x"5e",  x"f0",  x"97",  x"e5",  x"8a",  x"85",  x"8a",  x"e8", -- 10C8
         x"19",  x"e2",  x"d8",  x"d6",  x"85",  x"b4",  x"07",  x"bc", -- 10D0
         x"f6",  x"09",  x"90",  x"1a",  x"f1",  x"f1",  x"e5",  x"cd", -- 10D8
         x"55",  x"e5",  x"1b",  x"7d",  x"b4",  x"b7",  x"86",  x"46", -- 10E0
         x"2b",  x"4e",  x"e5",  x"b6",  x"67",  x"6e",  x"26",  x"46", -- 10E8
         x"aa",  x"d0",  x"2b",  x"56",  x"2e",  x"ae",  x"95",  x"b4", -- 10F0
         x"bf",  x"5d",  x"9b",  x"0e",  x"2b",  x"c3",  x"0c",  x"4d", -- 10F8
         x"ff",  x"bc",  x"39",  x"e7",  x"f5",  x"03",  x"e1",  x"91", -- 1100
         x"7e",  x"27",  x"c9",  x"85",  x"86",  x"1e",  x"1c",  x"da", -- 1108
         x"10",  x"86",  x"7b",  x"d1",  x"d1",  x"a7",  x"96",  x"cd", -- 1110
         x"16",  x"01",  x"d3",  x"15",  x"c2",  x"a8",  x"fc",  x"cd", -- 1118
         x"e9",  x"d2",  x"a6",  x"02",  x"21",  x"f2",  x"39",  x"62", -- 1120
         x"18",  x"6f",  x"ca",  x"6b",  x"ba",  x"e7",  x"6f",  x"2c", -- 1128
         x"a0",  x"00",  x"0a",  x"12",  x"03",  x"13",  x"18",  x"57", -- 1130
         x"f8",  x"3d",  x"3b",  x"df",  x"25",  x"e5",  x"99",  x"c0", -- 1138
         x"d5",  x"69",  x"1b",  x"4e",  x"28",  x"97",  x"70",  x"99", -- 1140
         x"47",  x"50",  x"09",  x"89",  x"e5",  x"90",  x"43",  x"ee", -- 1148
         x"61",  x"8a",  x"85",  x"89",  x"28",  x"14",  x"c0",  x"ea", -- 1150
         x"43",  x"c9",  x"01",  x"c0",  x"d0",  x"f0",  x"50",  x"fb", -- 1158
         x"d2",  x"af",  x"57",  x"a2",  x"80",  x"f2",  x"e9",  x"50", -- 1160
         x"0e",  x"30",  x"d3",  x"28",  x"55",  x"90",  x"da",  x"0c", -- 1168
         x"1a",  x"c9",  x"98",  x"b0",  x"80",  x"ca",  x"7f",  x"24", -- 1170
         x"d4",  x"7a",  x"6e",  x"73",  x"e0",  x"a9",  x"c0",  x"0a", -- 1178
         x"da",  x"d3",  x"af",  x"e3",  x"4f",  x"e5",  x"d7",  x"ef", -- 1180
         x"d8",  x"e0",  x"78",  x"11",  x"0e",  x"00",  x"f2",  x"2b", -- 1188
         x"ef",  x"1f",  x"c1",  x"e1",  x"e5",  x"2c",  x"cd",  x"45", -- 1190
         x"66",  x"68",  x"0e",  x"a2",  x"d8",  x"14",  x"d5",  x"56", -- 1198
         x"89",  x"76",  x"b3",  x"05",  x"18",  x"cf",  x"68",  x"2d", -- 11A0
         x"99",  x"1a",  x"39",  x"90",  x"18",  x"e3",  x"02",  x"7e", -- 11A8
         x"cd",  x"de",  x"d3",  x"04",  x"05",  x"98",  x"84",  x"c5", -- 11B0
         x"1e",  x"19",  x"ff",  x"fe",  x"29",  x"8b",  x"dc",  x"fa", -- 11B8
         x"af",  x"21",  x"92",  x"c3",  x"f1",  x"e3",  x"01",  x"61", -- 11C0
         x"cb",  x"33",  x"3d",  x"be",  x"3c",  x"6a",  x"d0",  x"cb", -- 11C8
         x"91",  x"05",  x"bb",  x"47",  x"d8",  x"43",  x"c9",  x"07", -- 11D0
         x"7f",  x"ca",  x"cf",  x"d4",  x"5f",  x"54",  x"22",  x"c3", -- 11D8
         x"06",  x"19",  x"46",  x"72",  x"e3",  x"eb",  x"75",  x"d2", -- 11E0
         x"b8",  x"67",  x"70",  x"c9",  x"eb",  x"ae",  x"31",  x"c2", -- 11E8
         x"55",  x"c5",  x"23",  x"80",  x"92",  x"4f",  x"ed",  x"78", -- 11F0
         x"60",  x"c3",  x"ad",  x"cd",  x"3e",  x"14",  x"d4",  x"81", -- 11F8
         x"07",  x"03",  x"4f",  x"7b",  x"ed",  x"79",  x"13",  x"b5", -- 1200
         x"0a",  x"f5",  x"c8",  x"bd",  x"f4",  x"99",  x"5e",  x"c1", -- 1208
         x"78",  x"19",  x"25",  x"ab",  x"a0",  x"28",  x"5f",  x"fa", -- 1210
         x"d3",  x"ba",  x"32",  x"0d",  x"17",  x"5e",  x"2b",  x"fd", -- 1218
         x"52",  x"80",  x"95",  x"61",  x"c9",  x"b7",  x"98",  x"8f", -- 1220
         x"53",  x"2e",  x"7b",  x"04",  x"e4",  x"c5",  x"1a",  x"18", -- 1228
         x"04",  x"b2",  x"cd",  x"6c",  x"c9",  x"d5",  x"a5",  x"38", -- 1230
         x"d1",  x"12",  x"b0",  x"12",  x"eb",  x"d4",  x"09",  x"7e", -- 1238
         x"c3",  x"b1",  x"d0",  x"f4",  x"16",  x"06",  x"e3",  x"88", -- 1240
         x"d3",  x"21",  x"28",  x"04",  x"d9",  x"9b",  x"ca",  x"18", -- 1248
         x"09",  x"04",  x"61",  x"21",  x"8b",  x"56",  x"fb",  x"78", -- 1250
         x"c9",  x"ff",  x"3a",  x"c3",  x"c5",  x"b7",  x"9d",  x"90", -- 1258
         x"d6",  x"90",  x"30",  x"0c",  x"15",  x"2f",  x"3c",  x"eb", -- 1260
         x"e0",  x"97",  x"97",  x"78",  x"1b",  x"fe",  x"19",  x"d0", -- 1268
         x"dc",  x"95",  x"03",  x"d7",  x"32",  x"67",  x"f1",  x"93", -- 1270
         x"19",  x"d5",  x"b4",  x"21",  x"96",  x"18",  x"f2",  x"ab", -- 1278
         x"f1",  x"00",  x"0a",  x"d5",  x"30",  x"4b",  x"23",  x"34", -- 1280
         x"28",  x"31",  x"63",  x"2e",  x"d8",  x"00",  x"3e",  x"d5", -- 1288
         x"18",  x"40",  x"af",  x"90",  x"47",  x"7e",  x"33",  x"9b", -- 1290
         x"5f",  x"67",  x"9a",  x"57",  x"03",  x"00",  x"99",  x"4f", -- 1298
         x"dc",  x"16",  x"d5",  x"68",  x"63",  x"af",  x"76",  x"47", -- 12A0
         x"a7",  x"20",  x"00",  x"16",  x"4a",  x"54",  x"65",  x"6f", -- 12A8
         x"78",  x"d6",  x"08",  x"0e",  x"fe",  x"e0",  x"20",  x"f0", -- 12B0
         x"86",  x"b0",  x"5d",  x"c9",  x"05",  x"29",  x"cb",  x"00", -- 12B8
         x"12",  x"cb",  x"11",  x"f2",  x"d4",  x"d4",  x"78",  x"5c", -- 12C0
         x"6a",  x"45",  x"cb",  x"08",  x"60",  x"21",  x"12",  x"86", -- 12C8
         x"77",  x"30",  x"e5",  x"c8",  x"78",  x"78",  x"08",  x"79", -- 12D0
         x"fc",  x"fd",  x"d4",  x"a0",  x"aa",  x"06",  x"e6",  x"80", -- 12D8
         x"a9",  x"4f",  x"c3",  x"76",  x"1c",  x"00",  x"c0",  x"14", -- 12E0
         x"c0",  x"0c",  x"c0",  x"0e",  x"80",  x"34",  x"02",  x"c0", -- 12E8
         x"c3",  x"53",  x"d6",  x"7e",  x"83",  x"94",  x"5b",  x"8a", -- 12F0
         x"5b",  x"89",  x"60",  x"4f",  x"b7",  x"e9",  x"c8",  x"e0", -- 12F8
         x"2f",  x"77",  x"36",  x"af",  x"6f",  x"71",  x"7d",  x"71", -- 1300
         x"7d",  x"dd",  x"70",  x"7d",  x"6f",  x"6f",  x"a0",  x"62", -- 1308
         x"a8",  x"b8",  x"43",  x"5a",  x"51",  x"c8",  x"ca",  x"18", -- 1310
         x"f5",  x"3a",  x"c6",  x"09",  x"f1",  x"cc",  x"c7",  x"79", -- 1318
         x"1f",  x"01",  x"4f",  x"cb",  x"1a",  x"cb",  x"1b",  x"cb", -- 1320
         x"18",  x"ab",  x"e6",  x"00",  x"00",  x"00",  x"81",  x"03", -- 1328
         x"aa",  x"56",  x"19",  x"80",  x"f1",  x"22",  x"00",  x"76", -- 1330
         x"80",  x"45",  x"aa",  x"38",  x"82",  x"cd",  x"97",  x"18", -- 1338
         x"d6",  x"b7",  x"ea",  x"b3",  x"f8",  x"73",  x"49",  x"01", -- 1340
         x"35",  x"80",  x"f4",  x"a6",  x"04",  x"90",  x"2a",  x"f5", -- 1348
         x"70",  x"af",  x"98",  x"6f",  x"e9",  x"80",  x"d1",  x"04", -- 1350
         x"cd",  x"f5",  x"d5",  x"21",  x"48",  x"c4",  x"a8",  x"66", -- 1358
         x"d4",  x"30",  x"21",  x"4c",  x"05",  x"ce",  x"d9",  x"01", -- 1360
         x"80",  x"fa",  x"1f",  x"3e",  x"1a",  x"c0",  x"fc",  x"0b", -- 1368
         x"d8",  x"32",  x"01",  x"31",  x"0c",  x"18",  x"72",  x"c7", -- 1370
         x"ad",  x"40",  x"30",  x"c8",  x"2e",  x"15",  x"58",  x"d6", -- 1378
         x"79",  x"32",  x"68",  x"f7",  x"a5",  x"22",  x"e5",  x"d2", -- 1380
         x"01",  x"81",  x"23",  x"50",  x"58",  x"21",  x"bc",  x"d4", -- 1388
         x"e5",  x"9b",  x"03",  x"d5",  x"e5",  x"04",  x"e5",  x"58", -- 1390
         x"d9",  x"88",  x"28",  x"80",  x"06",  x"2e",  x"08",  x"1f", -- 1398
         x"67",  x"79",  x"30",  x"0b",  x"d3",  x"f1",  x"21",  x"74", -- 13A0
         x"19",  x"92",  x"3a",  x"d3",  x"2b",  x"89",  x"80",  x"95", -- 13A8
         x"2d",  x"7c",  x"20",  x"65",  x"e4",  x"83",  x"41",  x"b1", -- 13B0
         x"85",  x"bc",  x"08",  x"e7",  x"01",  x"20",  x"84",  x"bb", -- 13B8
         x"65",  x"ec",  x"1a",  x"5a",  x"05",  x"ca",  x"4b",  x"c3", -- 13C0
         x"2e",  x"ff",  x"00",  x"5c",  x"34",  x"34",  x"2b",  x"7e", -- 13C8
         x"32",  x"14",  x"03",  x"a5",  x"04",  x"10",  x"87",  x"04", -- 13D0
         x"0c",  x"03",  x"41",  x"eb",  x"81",  x"a1",  x"57",  x"5f", -- 13D8
         x"32",  x"17",  x"ab",  x"d4",  x"c5",  x"b3",  x"f0",  x"0b", -- 13E0
         x"03",  x"de",  x"00",  x"15",  x"3f",  x"30",  x"07",  x"0d", -- 13E8
         x"b1",  x"9f",  x"37",  x"d2",  x"98",  x"d5",  x"79",  x"3c", -- 13F0
         x"3d",  x"01",  x"1f",  x"fa",  x"ec",  x"d4",  x"17",  x"cb", -- 13F8
         x"13",  x"63",  x"e1",  x"89",  x"e6",  x"10",  x"3a",  x"a8", -- 1400
         x"19",  x"17",  x"1d",  x"79",  x"b2",  x"39",  x"b3",  x"20", -- 1408
         x"f4",  x"a0",  x"eb",  x"02",  x"35",  x"e1",  x"20",  x"c7", -- 1410
         x"1e",  x"0a",  x"a3",  x"8f",  x"e8",  x"20",  x"ca",  x"7c", -- 1418
         x"d6",  x"7d",  x"a0",  x"11",  x"ae",  x"80",  x"47",  x"1f", -- 1420
         x"00",  x"a8",  x"78",  x"f2",  x"7b",  x"d6",  x"c6",  x"80", -- 1428
         x"77",  x"ad",  x"94",  x"a2",  x"e3",  x"7f",  x"77",  x"98", -- 1430
         x"40",  x"80",  x"2f",  x"0d",  x"e1",  x"b7",  x"e1",  x"f2", -- 1438
         x"ba",  x"18",  x"18",  x"8c",  x"2c",  x"eb",  x"95",  x"c1", -- 1440
         x"c6",  x"02",  x"38",  x"c7",  x"47",  x"43",  x"82",  x"59", -- 1448
         x"31",  x"8d",  x"16",  x"18",  x"bc",  x"a4",  x"79",  x"a9", -- 1450
         x"80",  x"e7",  x"03",  x"fe",  x"2f",  x"17",  x"9f",  x"c0", -- 1458
         x"59",  x"3c",  x"2f",  x"06",  x"88",  x"41",  x"bd",  x"46", -- 1460
         x"1d",  x"4f",  x"70",  x"88",  x"40",  x"23",  x"36",  x"80", -- 1468
         x"17",  x"c3",  x"28",  x"b9",  x"d4",  x"15",  x"f0",  x"21", -- 1470
         x"cf",  x"23",  x"7e",  x"ee",  x"59",  x"80",  x"4b",  x"93", -- 1478
         x"7c",  x"83",  x"7a",  x"0d",  x"8b",  x"dd",  x"99",  x"80", -- 1480
         x"49",  x"82",  x"11",  x"db",  x"0f",  x"18",  x"51",  x"03", -- 1488
         x"f6",  x"99",  x"ed",  x"53",  x"17",  x"ed",  x"43",  x"ed", -- 1490
         x"16",  x"df",  x"97",  x"8a",  x"09",  x"71",  x"82",  x"4e", -- 1498
         x"83",  x"23",  x"30",  x"c9",  x"11",  x"0b",  x"06",  x"04", -- 14A0
         x"1a",  x"77",  x"1a",  x"13",  x"23",  x"10",  x"ee",  x"58", -- 14A8
         x"42",  x"07",  x"37",  x"1f",  x"1a",  x"77",  x"3f",  x"1f", -- 14B0
         x"c6",  x"94",  x"77",  x"79",  x"09",  x"4f",  x"14",  x"1f", -- 14B8
         x"ae",  x"c9",  x"bf",  x"18",  x"5d",  x"21",  x"a0",  x"d6", -- 14C0
         x"51",  x"e5",  x"64",  x"79",  x"c8",  x"46",  x"22",  x"ae", -- 14C8
         x"79",  x"b0",  x"e0",  x"32",  x"d7",  x"1f",  x"a9",  x"c9", -- 14D0
         x"02",  x"23",  x"78",  x"be",  x"c0",  x"2b",  x"79",  x"94", -- 14D8
         x"03",  x"7a",  x"03",  x"7b",  x"18",  x"96",  x"c0",  x"e1", -- 14E0
         x"e2",  x"a8",  x"47",  x"b1",  x"70",  x"ae",  x"f0",  x"2a", -- 14E8
         x"c9",  x"a0",  x"de",  x"00",  x"ae",  x"67",  x"fc",  x"69", -- 14F0
         x"d7",  x"3e",  x"98",  x"90",  x"a4",  x"c8",  x"19",  x"7c", -- 14F8
         x"17",  x"dc",  x"ee",  x"e1",  x"ae",  x"49",  x"aa",  x"81", -- 1500
         x"23",  x"1b",  x"7a",  x"a3",  x"3c",  x"c0",  x"0b",  x"21", -- 1508
         x"8f",  x"8d",  x"fe",  x"98",  x"3a",  x"7e",  x"d0",  x"b0", -- 1510
         x"a7",  x"45",  x"d7",  x"36",  x"03",  x"98",  x"7b",  x"f5", -- 1518
         x"79",  x"17",  x"cd",  x"ca",  x"0e",  x"8a",  x"aa",  x"f9", -- 1520
         x"40",  x"78",  x"b1",  x"c8",  x"3e",  x"10",  x"29",  x"3d", -- 1528
         x"38",  x"06",  x"b6",  x"01",  x"eb",  x"30",  x"04",  x"09", -- 1530
         x"da",  x"0b",  x"d0",  x"ee",  x"de",  x"17",  x"fe",  x"00", -- 1538
         x"2d",  x"f5",  x"28",  x"05",  x"fe",  x"2b",  x"28",  x"01", -- 1540
         x"db",  x"8c",  x"ad",  x"16",  x"47",  x"67",  x"2f",  x"bf", -- 1548
         x"fc",  x"00",  x"38",  x"3d",  x"fe",  x"2e",  x"28",  x"16", -- 1550
         x"fe",  x"45",  x"2d",  x"20",  x"15",  x"a1",  x"8b",  x"4d", -- 1558
         x"ce",  x"12",  x"00",  x"4b",  x"14",  x"20",  x"07",  x"af", -- 1560
         x"93",  x"5f",  x"0c",  x"00",  x"0c",  x"28",  x"de",  x"e5", -- 1568
         x"7b",  x"90",  x"f4",  x"ed",  x"0d",  x"d7",  x"f2",  x"e4", -- 1570
         x"d7",  x"d2",  x"40",  x"e7",  x"d5",  x"f1",  x"3c",  x"20", -- 1578
         x"f2",  x"1a",  x"d1",  x"f1",  x"cc",  x"fb",  x"e2",  x"97", -- 1580
         x"c8",  x"cf",  x"0f",  x"82",  x"d6",  x"f0",  x"76",  x"a3", -- 1588
         x"0e",  x"57",  x"78",  x"89",  x"47",  x"c6",  x"56",  x"d5", -- 1590
         x"0d",  x"d6",  x"51",  x"30",  x"f4",  x"b3",  x"e1",  x"93", -- 1598
         x"28",  x"18",  x"a8",  x"a3",  x"ca",  x"cd",  x"a9",  x"9d", -- 15A0
         x"36",  x"c3",  x"85",  x"40",  x"7b",  x"07",  x"07",  x"83", -- 15A8
         x"07",  x"63",  x"86",  x"1a",  x"5f",  x"18",  x"a5",  x"d5", -- 15B0
         x"27",  x"0d",  x"d8",  x"35",  x"98",  x"59",  x"96",  x"9d", -- 15B8
         x"06",  x"98",  x"86",  x"62",  x"92",  x"c8",  x"65",  x"d1", -- 15C0
         x"11",  x"ea",  x"03",  x"8b",  x"96",  x"36",  x"57",  x"0c", -- 15C8
         x"42",  x"d8",  x"36",  x"2d",  x"8c",  x"80",  x"30",  x"ca", -- 15D0
         x"ef",  x"d8",  x"e5",  x"fc",  x"db",  x"60",  x"af",  x"5e", -- 15D8
         x"f5",  x"bf",  x"40",  x"43",  x"91",  x"11",  x"f8",  x"c0", -- 15E0
         x"a3",  x"18",  x"d7",  x"0d",  x"b7",  x"e2",  x"6e",  x"d8", -- 15E8
         x"d0",  x"18",  x"ee",  x"83",  x"12",  x"18",  x"ec",  x"05", -- 15F0
         x"85",  x"85",  x"1c",  x"cd",  x"5e",  x"d4",  x"3c",  x"05", -- 15F8
         x"f6",  x"23",  x"84",  x"01",  x"e0",  x"70",  x"f1",  x"81", -- 1600
         x"3c",  x"fa",  x"0c",  x"89",  x"d8",  x"fe",  x"08",  x"eb", -- 1608
         x"00",  x"3c",  x"47",  x"3e",  x"02",  x"3d",  x"3d",  x"00", -- 1610
         x"e1",  x"f5",  x"11",  x"08",  x"d9",  x"05",  x"20",  x"06", -- 1618
         x"28",  x"36",  x"2e",  x"52",  x"23",  x"05",  x"c5",  x"06", -- 1620
         x"cc",  x"f5",  x"d6",  x"86",  x"a4",  x"d5",  x"21",  x"e1", -- 1628
         x"06",  x"2f",  x"04",  x"8e",  x"e9",  x"9e",  x"c6",  x"7a", -- 1630
         x"9e",  x"9e",  x"c3",  x"79",  x"9e",  x"4f",  x"91",  x"a2", -- 1638
         x"30",  x"f0",  x"9d",  x"9c",  x"23",  x"5a",  x"46",  x"f0", -- 1640
         x"00",  x"70",  x"23",  x"c1",  x"0d",  x"20",  x"d2",  x"05", -- 1648
         x"34",  x"28",  x"0b",  x"bd",  x"38",  x"fe",  x"30",  x"bc", -- 1650
         x"c5",  x"97",  x"c4",  x"83",  x"35",  x"f1",  x"28",  x"1a", -- 1658
         x"36",  x"45",  x"44",  x"63",  x"2b",  x"81",  x"41",  x"9f", -- 1660
         x"bd",  x"e5",  x"00",  x"3d",  x"d6",  x"0a",  x"30",  x"fb", -- 1668
         x"c6",  x"3a",  x"23",  x"fd",  x"2c",  x"ed",  x"64",  x"71", -- 1670
         x"8b",  x"01",  x"05",  x"74",  x"94",  x"11",  x"f7",  x"23", -- 1678
         x"80",  x"a3",  x"e1",  x"e2",  x"65",  x"29",  x"d8",  x"e9", -- 1680
         x"bb",  x"80",  x"80",  x"a0",  x"86",  x"01",  x"10",  x"27", -- 1688
         x"64",  x"00",  x"9c",  x"00",  x"6e",  x"64",  x"0c",  x"0a", -- 1690
         x"02",  x"97",  x"eb",  x"9b",  x"e1",  x"d6",  x"e3",  x"e9", -- 1698
         x"43",  x"93",  x"70",  x"c3",  x"dd",  x"95",  x"b4",  x"40", -- 16A0
         x"78",  x"ca",  x"6d",  x"d9",  x"f2",  x"38",  x"29",  x"d9", -- 16A8
         x"b7",  x"bc",  x"73",  x"03",  x"d0",  x"d4",  x"ce",  x"61", -- 16B0
         x"79",  x"f6",  x"7f",  x"40",  x"9e",  x"f2",  x"29",  x"55", -- 16B8
         x"d9",  x"d9",  x"8d",  x"70",  x"d7",  x"23",  x"f5",  x"43", -- 16C0
         x"53",  x"e1",  x"7c",  x"1f",  x"a3",  x"fc",  x"af",  x"fc", -- 16C8
         x"03",  x"e3",  x"85",  x"dc",  x"1a",  x"d9",  x"0d",  x"f7", -- 16D0
         x"14",  x"1b",  x"59",  x"d5",  x"3f",  x"9a",  x"5b",  x"d5", -- 16D8
         x"85",  x"02",  x"38",  x"81",  x"11",  x"3b",  x"aa",  x"a9", -- 16E0
         x"0b",  x"e1",  x"01",  x"fe",  x"88",  x"d2",  x"76",  x"d6", -- 16E8
         x"5a",  x"37",  x"99",  x"e8",  x"fd",  x"da",  x"d6",  x"09", -- 16F0
         x"f5",  x"93",  x"ed",  x"61",  x"d5",  x"18",  x"91",  x"ac", -- 16F8
         x"db",  x"49",  x"6c",  x"09",  x"ca",  x"3b",  x"21",  x"ad", -- 1700
         x"7c",  x"52",  x"d9",  x"f9",  x"0c",  x"c1",  x"4a",  x"c3", -- 1708
         x"33",  x"08",  x"40",  x"00",  x"2e",  x"94",  x"74",  x"70", -- 1710
         x"4f",  x"2e",  x"77",  x"6e",  x"00",  x"02",  x"88",  x"7a", -- 1718
         x"e6",  x"a0",  x"2a",  x"7c",  x"50",  x"01",  x"aa",  x"aa", -- 1720
         x"7e",  x"ff",  x"ff",  x"7f",  x"7f",  x"40",  x"c0",  x"81", -- 1728
         x"b8",  x"81",  x"a0",  x"60",  x"11",  x"98",  x"d5",  x"d5", -- 1730
         x"91",  x"89",  x"35",  x"2e",  x"e1",  x"6f",  x"0e",  x"a3", -- 1738
         x"eb",  x"3f",  x"bb",  x"46",  x"50",  x"3d",  x"c8",  x"87", -- 1740
         x"0e",  x"f5",  x"18",  x"f5",  x"15",  x"95",  x"f2",  x"07", -- 1748
         x"e3",  x"30",  x"e1",  x"18",  x"dd",  x"a4",  x"e2",  x"00", -- 1750
         x"1b",  x"03",  x"fa",  x"5d",  x"da",  x"21",  x"3c",  x"03", -- 1758
         x"ec",  x"26",  x"0b",  x"c8",  x"86",  x"34",  x"e6",  x"07", -- 1760
         x"b0",  x"c4",  x"a4",  x"87",  x"87",  x"5d",  x"4f",  x"b4", -- 1768
         x"58",  x"a7",  x"03",  x"1a",  x"03",  x"3c",  x"e6",  x"03", -- 1770
         x"13",  x"0c",  x"fe",  x"01",  x"88",  x"32",  x"0a",  x"21", -- 1778
         x"60",  x"5d",  x"da",  x"1a",  x"86",  x"a6",  x"62",  x"7b", -- 1780
         x"0d",  x"59",  x"ee",  x"4f",  x"4f",  x"8a",  x"bd",  x"a4", -- 1788
         x"cd",  x"03",  x"21",  x"19",  x"b6",  x"80",  x"7e",  x"d6", -- 1790
         x"ab",  x"20",  x"04",  x"77",  x"0e",  x"0c",  x"15",  x"1c", -- 1798
         x"cd",  x"a3",  x"28",  x"50",  x"c3",  x"f7",  x"6d",  x"d6", -- 17A0
         x"e9",  x"4e",  x"01",  x"18",  x"a7",  x"80",  x"b1",  x"46", -- 17A8
         x"68",  x"99",  x"e9",  x"92",  x"00",  x"69",  x"10",  x"d1", -- 17B0
         x"75",  x"68",  x"21",  x"ba",  x"da",  x"ba",  x"3c",  x"88", -- 17B8
         x"12",  x"49",  x"83",  x"9a",  x"a3",  x"58",  x"8e",  x"58", -- 17C0
         x"f5",  x"99",  x"c8",  x"c0",  x"38",  x"f5",  x"6d",  x"3a", -- 17C8
         x"be",  x"21",  x"66",  x"6c",  x"db",  x"37",  x"35",  x"f2", -- 17D0
         x"a6",  x"09",  x"5e",  x"8c",  x"09",  x"b7",  x"f5",  x"f4", -- 17D8
         x"8a",  x"6f",  x"17",  x"39",  x"28",  x"f1",  x"d4",  x"09", -- 17E0
         x"c2",  x"da",  x"73",  x"c3",  x"b5",  x"ac",  x"3c",  x"49", -- 17E8
         x"f3",  x"00",  x"7f",  x"05",  x"ba",  x"d7",  x"1e",  x"86", -- 17F0
         x"03",  x"64",  x"26",  x"99",  x"87",  x"58",  x"34",  x"b6", -- 17F8
         x"00",  x"e0",  x"5d",  x"a5",  x"86",  x"6b",  x"da",  x"18", -- 1800
         x"83",  x"4f",  x"38",  x"76",  x"da",  x"b0",  x"9a",  x"df", -- 1808
         x"fd",  x"5b",  x"31",  x"f3",  x"ec",  x"64",  x"49",  x"fc", -- 1810
         x"91",  x"a9",  x"a8",  x"2c",  x"fb",  x"43",  x"81",  x"da", -- 1818
         x"09",  x"db",  x"e5",  x"21",  x"81",  x"51",  x"59",  x"75", -- 1820
         x"8c",  x"e8",  x"6f",  x"d4",  x"13",  x"55",  x"db",  x"8a", -- 1828
         x"50",  x"9e",  x"00",  x"c9",  x"09",  x"4a",  x"d7",  x"3b", -- 1830
         x"78",  x"02",  x"00",  x"6e",  x"84",  x"7b",  x"fe",  x"c1", -- 1838
         x"2f",  x"7c",  x"74",  x"00",  x"31",  x"9a",  x"7d",  x"84", -- 1840
         x"3d",  x"5a",  x"7d",  x"c8",  x"00",  x"7f",  x"91",  x"7e", -- 1848
         x"e4",  x"bb",  x"4c",  x"7e",  x"6c",  x"c5",  x"f1",  x"7f", -- 1850
         x"20",  x"e9",  x"85",  x"49",  x"db",  x"28",  x"03",  x"66", -- 1858
         x"e7",  x"37",  x"47",  x"6e",  x"db",  x"f1",  x"e9",  x"cc", -- 1860
         x"d3",  x"fe",  x"ae",  x"5c",  x"c0",  x"de",  x"ed",  x"88", -- 1868
         x"b0",  x"89",  x"0b",  x"fe",  x"94",  x"a6",  x"9c",  x"03", -- 1870
         x"47",  x"d2",  x"48",  x"c3",  x"d6",  x"07",  x"c3",  x"57", -- 1878
         x"da",  x"06",  x"b5",  x"d0",  x"00",  x"00",  x"b5",  x"6f", -- 1880
         x"eb",  x"18",  x"e0",  x"7b",  x"87",  x"a0",  x"00",  x"f6", -- 1888
         x"0d",  x"57",  x"1e",  x"33",  x"ef",  x"18",  x"be",  x"38", -- 1890
         x"e5",  x"36",  x"c9",  x"bf",  x"f0",  x"70",  x"f8",  x"b3", -- 1898
         x"cd",  x"03",  x"fe",  x"d2",  x"cd",  x"09",  x"d2",  x"2a", -- 18A0
         x"f6",  x"f0",  x"ed",  x"5b",  x"56",  x"03",  x"07",  x"af", -- 18A8
         x"ed",  x"52",  x"d1",  x"e3",  x"03",  x"9a",  x"14",  x"28", -- 18B0
         x"dd",  x"c8",  x"85",  x"e4",  x"dd",  x"47",  x"e1",  x"00", -- 18B8
         x"04",  x"12",  x"13",  x"2b",  x"7d",  x"b4",  x"20",  x"f6", -- 18C0
         x"b5",  x"0a",  x"5f",  x"28",  x"03",  x"57",  x"23",  x"38", -- 18C8
         x"44",  x"7f",  x"2a",  x"2b",  x"40",  x"0c",  x"90",  x"ae", -- 18D0
         x"1b",  x"7b",  x"b2",  x"fc",  x"1b",  x"33",  x"e8",  x"cc", -- 18D8
         x"f8",  x"dc",  x"38",  x"42",  x"20",  x"60",  x"2d",  x"26", -- 18E0
         x"77",  x"dd",  x"e3",  x"2b",  x"d5",  x"e9",  x"4c",  x"50", -- 18E8
         x"b8",  x"ce",  x"82",  x"05",  x"e1",  x"00",  x"42",  x"4b", -- 18F0
         x"03",  x"d1",  x"2b",  x"70",  x"2b",  x"71",  x"06",  x"2b", -- 18F8
         x"35",  x"03",  x"20",  x"fc",  x"ab",  x"b6",  x"76",  x"f0", -- 1900
         x"ca",  x"25",  x"fd",  x"dd",  x"d9",  x"69",  x"c0",  x"85", -- 1908
         x"18",  x"29",  x"00",  x"cd",  x"87",  x"dc",  x"e5",  x"e2", -- 1910
         x"7b",  x"db",  x"eb",  x"85",  x"ad",  x"7b",  x"5e",  x"e1", -- 1918
         x"80",  x"5e",  x"e1",  x"28",  x"c7",  x"cd",  x"1d",  x"de", -- 1920
         x"21",  x"00",  x"3f",  x"dc",  x"c3",  x"71",  x"c3",  x"42", -- 1928
         x"41",  x"44",  x"cc",  x"99",  x"ae",  x"28",  x"0c",  x"c6", -- 1930
         x"cd",  x"b0",  x"dc",  x"6c",  x"d7",  x"03",  x"2a",  x"1b", -- 1938
         x"1b",  x"c6",  x"03",  x"39",  x"01",  x"d1",  x"ff",  x"41", -- 1940
         x"14",  x"09",  x"44",  x"4d",  x"43",  x"6f",  x"a2",  x"3e", -- 1948
         x"67",  x"e5",  x"84",  x"33",  x"d2",  x"3e",  x"c3",  x"4e", -- 1950
         x"49",  x"91",  x"19",  x"2a",  x"21",  x"12",  x"6e",  x"d6", -- 1958
         x"c3",  x"0e",  x"8a",  x"c4",  x"1e",  x"26",  x"ae",  x"f6", -- 1960
         x"0a",  x"ac",  x"59",  x"cd",  x"01",  x"cc",  x"c8",  x"3b", -- 1968
         x"3e",  x"01",  x"32",  x"cc",  x"89",  x"d6",  x"06",  x"cf", -- 1970
         x"58",  x"05",  x"94",  x"8f",  x"60",  x"69",  x"eb",  x"d1", -- 1978
         x"19",  x"4e",  x"fa",  x"83",  x"09",  x"09",  x"23",  x"3a", -- 1980
         x"ae",  x"8f",  x"b0",  x"c9",  x"3e",  x"d4",  x"23",  x"00", -- 1988
         x"01",  x"3e",  x"d3",  x"f5",  x"3a",  x"5d",  x"03",  x"a7", -- 1990
         x"18",  x"3e",  x"00",  x"32",  x"05",  x"28",  x"04",  x"f1", -- 1998
         x"35",  x"c6",  x"04",  x"a8",  x"72",  x"be",  x"81",  x"3a", -- 19A0
         x"3c",  x"cd",  x"f1",  x"2e",  x"09",  x"3f",  x"d3",  x"78", -- 19A8
         x"21",  x"fe",  x"06",  x"38",  x"0d",  x"2b",  x"99",  x"00", -- 19B0
         x"10",  x"fb",  x"d5",  x"11",  x"82",  x"dc",  x"73",  x"23", -- 19B8
         x"0c",  x"72",  x"d1",  x"23",  x"f1",  x"9e",  x"6d",  x"01", -- 19C0
         x"eb",  x"80",  x"47",  x"79",  x"fe",  x"09",  x"38",  x"04", -- 19C8
         x"0d",  x"23",  x"0c",  x"18",  x"f7",  x"ed",  x"b0",  x"b7", -- 19D0
         x"bf",  x"ba",  x"74",  x"86",  x"ac",  x"dd",  x"32",  x"20", -- 19D8
         x"fa",  x"b9",  x"0b",  x"4f",  x"30",  x"01",  x"04",  x"81", -- 19E0
         x"13",  x"79",  x"c9",  x"5a",  x"1e",  x"07",  x"03",  x"cb", -- 19E8
         x"bc",  x"f8",  x"7d",  x"06",  x"3e",  x"13",  x"20",  x"02", -- 19F0
         x"02",  x"c6",  x"08",  x"32",  x"08",  x"03",  x"a0",  x"ec", -- 19F8
         x"f1",  x"c3",  x"2c",  x"d5",  x"dd",  x"19",  x"47",  x"cb", -- 1A00
         x"5a",  x"c7",  x"19",  x"12",  x"45",  x"19",  x"09",  x"b0", -- 1A08
         x"19",  x"c3",  x"d2",  x"a0",  x"fd",  x"67",  x"24",  x"d8", -- 1A10
         x"62",  x"80",  x"2a",  x"c0",  x"d4",  x"11",  x"ff",  x"30", -- 1A18
         x"fb",  x"19",  x"f7",  x"61",  x"11",  x"4f",  x"cd",  x"b5", -- 1A20
         x"dd",  x"e1",  x"9d",  x"9a",  x"0c",  x"33",  x"8e",  x"11", -- 1A28
         x"43",  x"cf",  x"0e",  x"f6",  x"df",  x"65",  x"84",  x"db", -- 1A30
         x"e2",  x"89",  x"50",  x"dd",  x"c1",  x"d0",  x"dd",  x"e6", -- 1A38
         x"87",  x"e5",  x"a7",  x"e0",  x"d8",  x"9a",  x"77",  x"34", -- 1A40
         x"77",  x"81",  x"f2",  x"60",  x"85",  x"f4",  x"ac",  x"1f", -- 1A48
         x"b1",  x"92",  x"c5",  x"d0",  x"1d",  x"3b",  x"c1",  x"79", -- 1A50
         x"cd",  x"ca",  x"72",  x"78",  x"eb",  x"04",  x"e3",  x"eb", -- 1A58
         x"95",  x"b0",  x"28",  x"b4",  x"56",  x"2b",  x"64",  x"5e", -- 1A60
         x"b8",  x"28",  x"28",  x"f3",  x"1a",  x"10",  x"13",  x"0b", -- 1A68
         x"fc",  x"fd",  x"23",  x"e5",  x"da",  x"1f",  x"0d",  x"1f", -- 1A70
         x"e1",  x"f1",  x"1f",  x"cf",  x"60",  x"1a",  x"aa",  x"f6", -- 1A78
         x"30",  x"c9",  x"3a",  x"a9",  x"db",  x"b9",  x"d4",  x"5f", -- 1A80
         x"46",  x"99",  x"23",  x"3e",  x"0c",  x"d1",  x"45",  x"57", -- 1A88
         x"14",  x"0f",  x"5f",  x"7a",  x"78",  x"7b",  x"e9",  x"d8", -- 1A90
         x"3c",  x"b3",  x"c3",  x"09",  x"0c",  x"ba",  x"0b",  x"b4", -- 1A98
         x"00",  x"7a",  x"18",  x"06",  x"d5",  x"29",  x"1e",  x"80", -- 1AA0
         x"0c",  x"cb",  x"e1",  x"19",  x"ef",  x"c8",  x"dd",  x"c5", -- 1AA8
         x"11",  x"42",  x"c4",  x"b1",  x"06",  x"7a",  x"b0",  x"aa", -- 1AB0
         x"31",  x"3e",  x"dc",  x"15",  x"1c",  x"10",  x"f8",  x"b0", -- 1AB8
         x"84",  x"e1",  x"3e",  x"f5",  x"a1",  x"df",  x"eb",  x"2b", -- 1AC0
         x"06",  x"8e",  x"2f",  x"47",  x"83",  x"ce",  x"d9",  x"45", -- 1AC8
         x"23",  x"20",  x"31",  x"21",  x"da",  x"30",  x"38",  x"ee", -- 1AD0
         x"79",  x"8b",  x"28",  x"50",  x"12",  x"2d",  x"87",  x"fe", -- 1AD8
         x"04",  x"c0",  x"07",  x"30",  x"16",  x"cb",  x"4e",  x"cb", -- 1AE0
         x"ce",  x"b1",  x"8e",  x"51",  x"3c",  x"27",  x"e1",  x"c3", -- 1AE8
         x"90",  x"89",  x"cb",  x"5e",  x"cb",  x"00",  x"de",  x"18", -- 1AF0
         x"ee",  x"cb",  x"6e",  x"cb",  x"ee",  x"18",  x"63",  x"e8", -- 1AF8
         x"e2",  x"da",  x"03",  x"39",  x"30",  x"a9",  x"39",  x"8b", -- 1B00
         x"63",  x"00",  x"3a",  x"10",  x"38",  x"14",  x"cb",  x"66", -- 1B08
         x"cb",  x"4c",  x"e6",  x"c9",  x"3c",  x"8a",  x"00",  x"c4", -- 1B10
         x"cb",  x"56",  x"cb",  x"d6",  x"18",  x"f0",  x"03",  x"cb", -- 1B18
         x"46",  x"cb",  x"c6",  x"18",  x"ea",  x"38",  x"f1",  x"03", -- 1B20
         x"8b",  x"78",  x"2a",  x"95",  x"23",  x"a0",  x"00",  x"01", -- 1B28
         x"61",  x"03",  x"c5",  x"ae",  x"c9",  x"31",  x"d7",  x"de", -- 1B30
         x"ae",  x"35",  x"fe",  x"22",  x"d6",  x"03",  x"b7",  x"28", -- 1B38
         x"1f",  x"f2",  x"a7",  x"de",  x"1d",  x"15",  x"9a",  x"c7", -- 1B40
         x"c1",  x"13",  x"80",  x"fa",  x"b7",  x"f2",  x"bb",  x"d3", -- 1B48
         x"70",  x"e4",  x"98",  x"1e",  x"d8",  x"b7",  x"ca",  x"80", -- 1B50
         x"3e",  x"20",  x"03",  x"18",  x"0c",  x"03",  x"02",  x"c4", -- 1B58
         x"fd",  x"56",  x"fc",  x"18",  x"09",  x"e1",  x"d0",  x"cb", -- 1B60
         x"28",  x"2a",  x"a5",  x"43",  x"af",  x"02",  x"e1",  x"77", -- 1B68
         x"7f",  x"cd",  x"a4",  x"c5",  x"9e",  x"8e",  x"ed",  x"94", -- 1B70
         x"9e",  x"74",  x"8a",  x"80",  x"fe",  x"0a",  x"20",  x"05", -- 1B78
         x"cd",  x"2b",  x"12",  x"df",  x"db",  x"cc",  x"0f",  x"df", -- 1B80
         x"c0",  x"cf",  x"27",  x"df",  x"9b",  x"00",  x"32",  x"df", -- 1B88
         x"18",  x"e7",  x"fe",  x"0d",  x"14",  x"c0",  x"3e",  x"09", -- 1B90
         x"30",  x"23",  x"6a",  x"7e",  x"49",  x"f6",  x"d1",  x"b6", -- 1B98
         x"20",  x"a1",  x"1b",  x"30",  x"c3",  x"d4",  x"06",  x"fe", -- 1BA0
         x"ba",  x"07",  x"02",  x"a7",  x"2a",  x"b6",  x"2f",  x"37", -- 1BA8
         x"e8",  x"19",  x"08",  x"28",  x"44",  x"c8",  x"80",  x"28", -- 1BB0
         x"2a",  x"fe",  x"1f",  x"28",  x"47",  x"fe",  x"00",  x"19", -- 1BB8
         x"ca",  x"c5",  x"df",  x"fe",  x"18",  x"ca",  x"cf",  x"c6", -- 1BC0
         x"04",  x"02",  x"ca",  x"db",  x"04",  x"1a",  x"07",  x"28", -- 1BC8
         x"48",  x"fe",  x"0b",  x"c8",  x"5a",  x"bc",  x"02",  x"01", -- 1BD0
         x"02",  x"f8",  x"0a",  x"05",  x"3f",  x"4a",  x"25",  x"c9", -- 1BD8
         x"77",  x"4f",  x"dc",  x"9e",  x"ab",  x"03",  x"a3",  x"e5", -- 1BE0
         x"3a",  x"28",  x"07",  x"7e",  x"84",  x"0a",  x"d2",  x"03", -- 1BE8
         x"a2",  x"c6",  x"60",  x"f0",  x"15",  x"6e",  x"18",  x"df", -- 1BF0
         x"e5",  x"23",  x"a0",  x"9a",  x"f4",  x"fb",  x"c6",  x"d1", -- 1BF8
         x"73",  x"af",  x"cb",  x"e3",  x"2d",  x"17",  x"78",  x"20", -- 1C00
         x"f7",  x"6b",  x"ec",  x"0e",  x"b0",  x"25",  x"34",  x"2a", -- 1C08
         x"20",  x"0c",  x"15",  x"af",  x"11",  x"33",  x"3b",  x"67", -- 1C10
         x"d1",  x"e2",  x"f9",  x"c4",  x"02",  x"0b",  x"7e",  x"0c", -- 1C18
         x"28",  x"4b",  x"20",  x"4b",  x"c9",  x"4a",  x"4c",  x"c1", -- 1C20
         x"b2",  x"89",  x"bc",  x"00",  x"18",  x"90",  x"cd",  x"c5", -- 1C28
         x"ff",  x"58",  x"09",  x"bc",  x"eb",  x"6f",  x"f2",  x"45", -- 1C30
         x"e1",  x"f6",  x"61",  x"10",  x"fe",  x"00",  x"c9",  x"1e", -- 1C38
         x"ff",  x"c3",  x"0e",  x"25",  x"e0",  x"ff",  x"00",  x"80", -- 1C40
         x"00",  x"40",  x"d5",  x"00",  x"2e",  x"08",  x"e5",  x"3e", -- 1C48
         x"01",  x"cd",  x"04",  x"e4",  x"00",  x"7c",  x"3c",  x"28", -- 1C50
         x"0f",  x"7d",  x"cd",  x"59",  x"f3",  x"50",  x"7c",  x"03", -- 1C58
         x"7a",  x"cd",  x"76",  x"00",  x"f3",  x"cd",  x"6b",  x"f3", -- 1C60
         x"e1",  x"7d",  x"c6",  x"04",  x"14",  x"6f",  x"30",  x"e0", -- 1C68
         x"09",  x"d1",  x"00",  x"c9",  x"d5",  x"cd",  x"ee",  x"f1", -- 1C70
         x"43",  x"41",  x"4f",  x"00",  x"53",  x"00",  x"3e",  x"45", -- 1C78
         x"cd",  x"29",  x"e3",  x"db",  x"00",  x"88",  x"0f",  x"38", -- 1C80
         x"05",  x"cd",  x"ec",  x"c0",  x"18",  x"0a",  x"03",  x"cd", -- 1C88
         x"e2",  x"c0",  x"19",  x"00",  x"52",  x"4f",  x"4d",  x"43", -- 1C90
         x"20",  x"00",  x"dd",  x"7e",  x"13",  x"04",  x"cb",  x"3f", -- 1C98
         x"89",  x"01",  x"2f",  x"e6",  x"33",  x"08",  x"28",  x"5f", -- 1CA0
         x"07",  x"a0",  x"29",  x"da",  x"c0",  x"3e",  x"30",  x"a1", -- 1CA8
         x"15",  x"cb",  x"4b",  x"20",  x"18",  x"13",  x"34",  x"a0", -- 1CB0
         x"13",  x"dd",  x"cb",  x"04",  x"46",  x"8c",  x"15",  x"a5", -- 1CB8
         x"56",  x"38",  x"a7",  x"53",  x"01",  x"51",  x"2c",  x"c6", -- 1CC0
         x"2e",  x"50",  x"89",  x"cb",  x"44",  x"6f",  x"d2",  x"26", -- 1CC8
         x"1d",  x"5f",  x"83",  x"27",  x"42",  x"49",  x"4c",  x"44", -- 1CD0
         x"2a",  x"31",  x"cb",  x"53",  x"5c",  x"28",  x"01",  x"3c", -- 1CD8
         x"52",  x"24",  x"05",  x"b1",  x"80",  x"96",  x"41",  x"4d", -- 1CE0
         x"00",  x"b0",  x"07",  x"20",  x"4f",  x"4e",  x"0d",  x"4c", -- 1CE8
         x"0a",  x"09",  x"46",  x"58",  x"46",  x"0a",  x"21",  x"00", -- 1CF0
         x"b9",  x"01",  x"01",  x"f0",  x"0c",  x"0c",  x"79",  x"cd", -- 1CF8
         x"eb",  x"82",  x"12",  x"3a",  x"00",  x"cd",  x"cf",  x"f6", -- 1D00
         x"80",  x"32",  x"10",  x"f0",  x"c9",  x"af",  x"3e",  x"ff", -- 1D08
         x"00",  x"5f",  x"57",  x"3c",  x"13",  x"13",  x"ed",  x"52", -- 1D10
         x"f2",  x"00",  x"13",  x"c1",  x"c9",  x"06",  x"00",  x"1e", -- 1D18
         x"09",  x"7a",  x"00",  x"1f",  x"1d",  x"c8",  x"57",  x"78", -- 1D20
         x"30",  x"01",  x"81",  x"00",  x"1f",  x"47",  x"18",  x"f3", -- 1D28
         x"f5",  x"fe",  x"0a",  x"30",  x"00",  x"2e",  x"7a",  x"a7", -- 1D30
         x"28",  x"2a",  x"84",  x"38",  x"27",  x"06",  x"fe",  x"21", -- 1D38
         x"30",  x"23",  x"7b",  x"0a",  x"1f",  x"00",  x"85",  x"38", -- 1D40
         x"1c",  x"fe",  x"29",  x"30",  x"18",  x"f1",  x"00",  x"d5", -- 1D48
         x"e5",  x"cd",  x"bb",  x"f6",  x"e1",  x"d1",  x"22",  x"06", -- 1D50
         x"9c",  x"b7",  x"ed",  x"53",  x"9e",  x"03",  x"43",  x"00", -- 1D58
         x"a0",  x"b7",  x"32",  x"9b",  x"b7",  x"a7",  x"c9",  x"f1", -- 1D60
         x"03",  x"37",  x"c9",  x"3e",  x"1f",  x"a5",  x"17",  x"00", -- 1D68
         x"00",  x"6f",  x"3a",  x"81",  x"b7",  x"fe",  x"02",  x"7b", -- 1D70
         x"30",  x"00",  x"03",  x"3a",  x"a3",  x"b7",  x"e6",  x"07", -- 1D78
         x"b5",  x"32",  x"de",  x"05",  x"c9",  x"46",  x"27",  x"5b", -- 1D80
         x"05",  x"88",  x"b7",  x"d9",  x"2a",  x"82",  x"0c",  x"07", -- 1D88
         x"86",  x"b7",  x"af",  x"75",  x"30",  x"07",  x"18",  x"19", -- 1D90
         x"eb",  x"d9",  x"01",  x"18",  x"f4",  x"d9",  x"53",  x"d5", -- 1D98
         x"0c",  x"06",  x"0c",  x"00",  x"f6",  x"01",  x"18",  x"f6", -- 1DA0
         x"e5",  x"d9",  x"c1",  x"e5",  x"0c",  x"ed",  x"42",  x"e1", -- 1DA8
         x"c5",  x"3a",  x"e3",  x"f6",  x"0c",  x"02",  x"e5",  x"44", -- 1DB0
         x"4d",  x"0e",  x"d1",  x"60",  x"00",  x"69",  x"cb",  x"3c", -- 1DB8
         x"cb",  x"1d",  x"d9",  x"e1",  x"eb",  x"05",  x"cd",  x"e8", -- 1DC0
         x"f7",  x"d9",  x"a7",  x"00",  x"2a",  x"01",  x"09",  x"d9", -- 1DC8
         x"cb",  x"4f",  x"20",  x"04",  x"00",  x"23",  x"30",  x"0b", -- 1DD0
         x"a7",  x"cb",  x"47",  x"13",  x"28",  x"18",  x"02",  x"1b", -- 1DD8
         x"1b",  x"12",  x"23",  x"08",  x"78",  x"00",  x"b1",  x"c8", -- 1DE0
         x"0b",  x"08",  x"18",  x"db",  x"e5",  x"d5",  x"07",  x"c5", -- 1DE8
         x"2a",  x"d3",  x"b7",  x"7d",  x"75",  x"73",  x"34",  x"80", -- 1DF0
         x"03",  x"c6",  x"f8",  x"4f",  x"06",  x"fd",  x"3a",  x"d5", -- 1DF8
         x"00",  x"b7",  x"2f",  x"67",  x"0a",  x"cd",  x"4e",  x"e0", -- 1E00
         x"38",  x"02",  x"16",  x"47",  x"4e",  x"2f",  x"a1",  x"77", -- 1E08
         x"c4",  x"cf",  x"ee",  x"02",  x"06",  x"f3",  x"d3",  x"84", -- 1E10
         x"56",  x"7b",  x"03",  x"fb",  x"1b",  x"78",  x"a1",  x"7a", -- 1E18
         x"6a",  x"e1",  x"b6",  x"10",  x"54",  x"f3",  x"e5",  x"41", -- 1E20
         x"0a",  x"cd",  x"4a",  x"f6",  x"23",  x"99",  x"30",  x"10", -- 1E28
         x"f7",  x"e1",  x"41",  x"04",  x"3e",  x"09",  x"cd",  x"1d", -- 1E30
         x"f2",  x"86",  x"0f",  x"2a",  x"f6",  x"0f",  x"c9",  x"03", -- 1E38
         x"fe",  x"03",  x"30",  x"08",  x"0e",  x"08",  x"da",  x"00", -- 1E40
         x"30",  x"02",  x"1e",  x"04",  x"cc",  x"a5",  x"23",  x"c2", -- 1E48
         x"a1",  x"c9",  x"01",  x"cd",  x"de",  x"e3",  x"38",  x"06", -- 1E50
         x"1d",  x"20",  x"8c",  x"24",  x"17",  x"f2",  x"d1",  x"1e", -- 1E58
         x"c8",  x"fe",  x"01",  x"13",  x"20",  x"e6",  x"18",  x"02", -- 1E60
         x"0e",  x"01",  x"43",  x"1c",  x"3e",  x"05",  x"32",  x"98", -- 1E68
         x"13",  x"cd",  x"34",  x"50",  x"01",  x"cd",  x"92",  x"f3", -- 1E70
         x"7e",  x"e1",  x"38",  x"51",  x"88",  x"c0",  x"ea",  x"2a", -- 1E78
         x"97",  x"48",  x"b7",  x"0d",  x"a7",  x"61",  x"23",  x"10", -- 1E80
         x"28",  x"04",  x"cd",  x"62",  x"8d",  x"57",  x"1a",  x"fe", -- 1E88
         x"2e",  x"33",  x"2c",  x"90",  x"e5",  x"13",  x"1a",  x"13", -- 1E90
         x"00",  x"18",  x"ef",  x"fe",  x"3a",  x"20",  x"03",  x"2b", -- 1E98
         x"18",  x"02",  x"c4",  x"fe",  x"2f",  x"20",  x"0b",  x"13", -- 1EA0
         x"8a",  x"26",  x"38",  x"1e",  x"2f",  x"02",  x"18",  x"b5", -- 1EA8
         x"fe",  x"27",  x"20",  x"0e",  x"b6",  x"1e",  x"3e",  x"ab", -- 1EB0
         x"09",  x"28",  x"19",  x"cf",  x"77",  x"23",  x"9b",  x"60", -- 1EB8
         x"0a",  x"a0",  x"fe",  x"20",  x"28",  x"b5",  x"03",  x"cd", -- 1EC0
         x"61",  x"f3",  x"18",  x"97",  x"21",  x"ea",  x"15",  x"7e", -- 1EC8
         x"00",  x"96",  x"24",  x"06",  x"08",  x"00",  x"cd",  x"b1", -- 1ED0
         x"c3",  x"38",  x"56",  x"21",  x"e2",  x"f9",  x"00",  x"22", -- 1ED8
         x"99",  x"b7",  x"11",  x"06",  x"fa",  x"21",  x"e1",  x"06", -- 1EE0
         x"b7",  x"cb",  x"4e",  x"20",  x"06",  x"a0",  x"4d",  x"be", -- 1EE8
         x"42",  x"04",  x"80",  x"05",  x"c4",  x"b7",  x"c3",  x"8f", -- 1EF0
         x"c3",  x"23",  x"46",  x"b3",  x"23",  x"32",  x"23",  x"7d", -- 1EF8
         x"0a",  x"3d",  x"20",  x"0a",  x"3a",  x"20",  x"33",  x"97", -- 1F00
         x"32",  x"04",  x"18",  x"0b",  x"0c",  x"5a",  x"1f",  x"0c", -- 1F08
         x"d7",  x"ba",  x"0c",  x"1a",  x"3a",  x"f5",  x"1d",  x"11", -- 1F10
         x"0f",  x"b0",  x"38",  x"11",  x"10",  x"1a",  x"cb",  x"8f", -- 1F18
         x"12",  x"0d",  x"18",  x"10",  x"18",  x"72",  x"11",  x"fb", -- 1F20
         x"72",  x"44",  x"16",  x"11",  x"cf",  x"12",  x"df",  x"4c", -- 1F28
         x"04",  x"2b",  x"38",  x"3c",  x"c0",  x"c9",  x"28",  x"1c", -- 1F30
         x"1a",  x"3d",  x"28",  x"0a",  x"1d",  x"51",  x"c5",  x"41", -- 1F38
         x"c7",  x"18",  x"05",  x"bf",  x"06",  x"87",  x"48",  x"28", -- 1F40
         x"87",  x"0f",  x"2f",  x"88",  x"0b",  x"28",  x"14",  x"05", -- 1F48
         x"20",  x"15",  x"71",  x"cb",  x"4a",  x"27",  x"01",  x"4f", -- 1F50
         x"a1",  x"21",  x"e6",  x"0f",  x"b1",  x"40",  x"22",  x"cd", -- 1F58
         x"d4",  x"fa",  x"3e",  x"0c",  x"00",  x"c5",  x"81",  x"06", -- 1F60
         x"02",  x"4f",  x"2a",  x"e2",  x"b7",  x"01",  x"f3",  x"ed", -- 1F68
         x"b3",  x"c1",  x"3a",  x"e4",  x"b7",  x"83",  x"79",  x"47", -- 1F70
         x"3e",  x"0a",  x"81",  x"4f",  x"0c",  x"18",  x"fb",  x"c9", -- 1F78
         x"c3",  x"dd",  x"00",  x"16",  x"3c",  x"0e",  x"80",  x"ed", -- 1F80
         x"78",  x"fe",  x"0a",  x"ee",  x"28",  x"09",  x"04",  x"00", -- 1F88
         x"19",  x"15",  x"20",  x"f3",  x"e0",  x"82",  x"e5",  x"68", -- 1F90
         x"3e",  x"02",  x"16",  x"d9",  x"c3",  x"e1",  x"ac",  x"0a", -- 1F98
         x"d5",  x"6c",  x"47",  x"c2",  x"0c",  x"25",  x"c4",  x"2a", -- 1FA0
         x"b9",  x"d0",  x"c0",  x"b6",  x"20",  x"1a",  x"11",  x"03", -- 1FA8
         x"fa",  x"c0",  x"3f",  x"28",  x"05",  x"21",  x"a3",  x"fb", -- 1FB0
         x"18",  x"1a",  x"18",  x"21",  x"a2",  x"04",  x"19",  x"c2", -- 1FB8
         x"c3",  x"cb",  x"08",  x"14",  x"3d",  x"90",  x"13",  x"a0", -- 1FC0
         x"fb",  x"1c",  x"58",  x"06",  x"c4",  x"58",  x"8f",  x"ee", -- 1FC8
         x"18",  x"22",  x"34",  x"88",  x"f0",  x"1b",  x"5b",  x"01", -- 1FD0
         x"31",  x"31",  x"61",  x"5b",  x"30",  x"31",  x"65",  x"80", -- 1FD8
         x"08",  x"37",  x"38",  x"71",  x"4b",  x"40",  x"02",  x"c5", -- 1FE0
         x"5b",  x"f5",  x"55",  x"7f",  x"f7",  x"40",  x"2a",  x"cb", -- 1FE8
         x"b7",  x"06",  x"c4",  x"f8",  x"28",  x"7e",  x"03",  x"23", -- 1FF0
         x"a7",  x"20",  x"02",  x"3e",  x"20",  x"ef",  x"15",  x"30", -- 1FF8
         x"30",  x"05",  x"cd",  x"46",  x"0d",  x"20",  x"ed",  x"3e", -- 2000
         x"18",  x"0d",  x"cd",  x"38",  x"ba",  x"28",  x"0a",  x"04", -- 2008
         x"10",  x"df",  x"00",  x"f1",  x"c3",  x"34",  x"f2",  x"e6", -- 2010
         x"f0",  x"28",  x"15",  x"0c",  x"fe",  x"10",  x"28",  x"5c", -- 2018
         x"23",  x"ca",  x"32",  x"06",  x"c5",  x"fe",  x"30",  x"ca", -- 2020
         x"b7",  x"04",  x"50",  x"00",  x"ca",  x"fa",  x"c5",  x"18", -- 2028
         x"e3",  x"26",  x"00",  x"e5",  x"0c",  x"21",  x"16",  x"c6", -- 2030
         x"06",  x"29",  x"0e",  x"c6",  x"02",  x"e1",  x"cd",  x"8f", -- 2038
         x"c4",  x"30",  x"f1",  x"97",  x"39",  x"51",  x"39",  x"80", -- 2040
         x"04",  x"c3",  x"54",  x"c4",  x"2e",  x"00",  x"01",  x"08", -- 2048
         x"c5",  x"20",  x"11",  x"00",  x"b7",  x"21",  x"93",  x"ed", -- 2050
         x"b0",  x"9e",  x"d6",  x"c1",  x"5b",  x"a9",  x"60",  x"79", -- 2058
         x"16",  x"17",  x"23",  x"10",  x"fa",  x"ac",  x"20",  x"67", -- 2060
         x"ef",  x"e1",  x"00",  x"2c",  x"3e",  x"28",  x"bd",  x"20", -- 2068
         x"da",  x"7c",  x"c6",  x"16",  x"08",  x"67",  x"c9",  x"4a", -- 2070
         x"20",  x"9b",  x"4a",  x"38",  x"26",  x"06",  x"04",  x"37", -- 2078
         x"18",  x"7e",  x"12",  x"13",  x"01",  x"2c",  x"10",  x"f8", -- 2080
         x"8f",  x"3d",  x"91",  x"40",  x"ec",  x"2b",  x"40",  x"d2", -- 2088
         x"40",  x"1b",  x"04",  x"67",  x"30",  x"c4",  x"8a",  x"82", -- 2090
         x"e5",  x"c5",  x"31",  x"db",  x"e8",  x"6b",  x"61",  x"c1", -- 2098
         x"f7",  x"9d",  x"0b",  x"2e",  x"80",  x"0a",  x"1b",  x"44", -- 20A0
         x"1a",  x"a5",  x"c7",  x"80",  x"37",  x"cb",  x"10",  x"13", -- 20A8
         x"3e",  x"06",  x"bb",  x"c5",  x"df",  x"a7",  x"a8",  x"08", -- 20B0
         x"78",  x"3a",  x"cb",  x"0d",  x"0a",  x"cb",  x"7d",  x"28", -- 20B8
         x"e1",  x"25",  x"37",  x"21",  x"2a",  x"72",  x"0e",  x"72", -- 20C0
         x"bb",  x"04",  x"2a",  x"5c",  x"2c",  x"0f",  x"0e",  x"06", -- 20C8
         x"cd",  x"00",  x"44",  x"b4",  x"29",  x"19",  x"57",  x"ef", -- 20D0
         x"32",  x"84",  x"67",  x"87",  x"8b",  x"49",  x"3f",  x"25", -- 20D8
         x"30",  x"92",  x"ea",  x"da",  x"d4",  x"25",  x"04",  x"25", -- 20E0
         x"af",  x"a0",  x"99",  x"9c",  x"29",  x"eb",  x"c3",  x"23", -- 20E8
         x"82",  x"c4",  x"03",  x"b0",  x"9b",  x"04",  x"f7",  x"2e", -- 20F0
         x"82",  x"0d",  x"78",  x"be",  x"ec",  x"bf",  x"26",  x"84", -- 20F8
         x"05",  x"df",  x"82",  x"84",  x"38",  x"60",  x"84",  x"50", -- 2100
         x"55",  x"84",  x"39",  x"0e",  x"8a",  x"60",  x"7d",  x"81", -- 2108
         x"8f",  x"94",  x"57",  x"f2",  x"24",  x"ec",  x"00",  x"80", -- 2110
         x"27",  x"21",  x"f2",  x"2c",  x"90",  x"d7",  x"fa",  x"20", -- 2118
         x"96",  x"7c",  x"65",  x"24",  x"ee",  x"58",  x"7c",  x"bd", -- 2120
         x"b4",  x"46",  x"23",  x"09",  x"41",  x"88",  x"56",  x"13", -- 2128
         x"d8",  x"54",  x"64",  x"10",  x"00",  x"f9",  x"c9",  x"0d", -- 2130
         x"09",  x"1b",  x"4a",  x"18",  x"1b",  x"09",  x"2a",  x"05", -- 2138
         x"40",  x"01",  x"db",  x"09",  x"80",  x"d2",  x"ca",  x"91", -- 2140
         x"60",  x"31",  x"32",  x"60",  x"1b",  x"4b",  x"e2",  x"17", -- 2148
         x"f9",  x"0d",  x"1b",  x"6a",  x"25",  x"16",  x"d0",  x"db", -- 2150
         x"03",  x"38",  x"38",  x"29",  x"21",  x"d1",  x"b5",  x"d6", -- 2158
         x"69",  x"da",  x"ae",  x"a1",  x"e5",  x"3a",  x"e8",  x"93", -- 2160
         x"82",  x"46",  x"d5",  x"5c",  x"b0",  x"f5",  x"cc",  x"52", -- 2168
         x"47",  x"f3",  x"33",  x"d6",  x"07",  x"88",  x"28",  x"03", -- 2170
         x"19",  x"c8",  x"78",  x"32",  x"17",  x"18",  x"06",  x"28", -- 2178
         x"24",  x"11",  x"78",  x"fa",  x"17",  x"01",  x"98",  x"fa", -- 2180
         x"28",  x"c2",  x"c3",  x"0a",  x"d3",  x"87",  x"be",  x"96", -- 2188
         x"c1",  x"1c",  x"08",  x"b4",  x"97",  x"d8",  x"09",  x"c7", -- 2190
         x"a2",  x"a2",  x"e1",  x"15",  x"94",  x"e5",  x"2a",  x"94", -- 2198
         x"a2",  x"e7",  x"d5",  x"94",  x"21",  x"b0",  x"3d",  x"22", -- 21A0
         x"28",  x"0e",  x"0d",  x"21",  x"01",  x"74",  x"c7",  x"22", -- 21A8
         x"1e",  x"06",  x"00",  x"0b",  x"0e",  x"0b",  x"18",  x"e6", -- 21B0
         x"21",  x"f0",  x"c6",  x"05",  x"11",  x"01",  x"a8",  x"01", -- 21B8
         x"11",  x"14",  x"da",  x"8e",  x"86",  x"d8",  x"f0",  x"e5", -- 21C0
         x"32",  x"00",  x"0d",  x"a8",  x"c9",  x"47",  x"5b",  x"b4", -- 21C8
         x"5b",  x"03",  x"da",  x"8d",  x"6a",  x"47",  x"2e",  x"f1", -- 21D0
         x"04",  x"44",  x"03",  x"e1",  x"82",  x"08",  x"02",  x"e2", -- 21D8
         x"14",  x"c7",  x"0a",  x"ea",  x"11",  x"18",  x"e6",  x"5a", -- 21E0
         x"b4",  x"a9",  x"02",  x"e5",  x"c0",  x"d8",  x"7e",  x"b7", -- 21E8
         x"c8",  x"23",  x"03",  x"2c",  x"7e",  x"02",  x"03",  x"2e", -- 21F0
         x"81",  x"00",  x"34",  x"7e",  x"c6",  x"f5",  x"30",  x"e9", -- 21F8
         x"c9",  x"5a",  x"72",  x"57",  x"c7",  x"cb",  x"1e",  x"5b", -- 2200
         x"28",  x"29",  x"a9",  x"00",  x"07",  x"ce",  x"3e",  x"d5", -- 2208
         x"be",  x"d5",  x"11",  x"38",  x"a0",  x"00",  x"9a",  x"d8", -- 2210
         x"5f",  x"05",  x"a6",  x"14",  x"d8",  x"b7",  x"b1",  x"45", -- 2218
         x"01",  x"0b",  x"00",  x"6a",  x"eb",  x"d1",  x"72",  x"3e", -- 2220
         x"74",  x"cd",  x"9c",  x"72",  x"c8",  x"b7",  x"cb",  x"74", -- 2228
         x"9b",  x"df",  x"da",  x"06",  x"b7",  x"72",  x"cb",  x"73", -- 2230
         x"20",  x"81",  x"2c",  x"dc",  x"ae",  x"0a",  x"20",  x"ea", -- 2238
         x"36",  x"df",  x"fb",  x"89",  x"00",  x"81",  x"c8",  x"cd", -- 2240
         x"95",  x"14",  x"c8",  x"18",  x"df",  x"0d",  x"8e",  x"38", -- 2248
         x"cd",  x"1c",  x"f8",  x"48",  x"88",  x"0e",  x"d0",  x"bd", -- 2250
         x"1c",  x"a5",  x"aa",  x"10",  x"b3",  x"d6",  x"21",  x"31", -- 2258
         x"ed",  x"4b",  x"51",  x"cd",  x"d9",  x"e4",  x"c9",  x"cd", -- 2260
         x"ff",  x"f5",  x"41",  x"18",  x"ae",  x"d1",  x"18",  x"de", -- 2268
         x"26",  x"7b",  x"4a",  x"ed",  x"a6",  x"7f",  x"66",  x"c8", -- 2270
         x"03",  x"dd",  x"77",  x"03",  x"39",  x"03",  x"8e",  x"e5", -- 2278
         x"e1",  x"da",  x"71",  x"c8",  x"b1",  x"a0",  x"02",  x"fe", -- 2280
         x"01",  x"c2",  x"ac",  x"07",  x"27",  x"be",  x"dd",  x"50", -- 2288
         x"34",  x"8e",  x"6c",  x"a0",  x"0b",  x"e5",  x"bf",  x"d5", -- 2290
         x"dd",  x"8a",  x"1e",  x"10",  x"ee",  x"c6",  x"98",  x"05", -- 2298
         x"12",  x"1a",  x"d6",  x"04",  x"98",  x"de",  x"12",  x"32", -- 22A0
         x"5e",  x"52",  x"03",  x"12",  x"f6",  x"ce",  x"da",  x"b4", -- 22A8
         x"a1",  x"be",  x"28",  x"b0",  x"20",  x"fe",  x"23",  x"13", -- 22B0
         x"10",  x"55",  x"f1",  x"af",  x"50",  x"0a",  x"7e",  x"c2", -- 22B8
         x"7b",  x"05",  x"f8",  x"eb",  x"3e",  x"75",  x"56",  x"02", -- 22C0
         x"bb",  x"7a",  x"70",  x"bc",  x"b0",  x"b7",  x"c1",  x"72", -- 22C8
         x"cd",  x"91",  x"e5",  x"38",  x"39",  x"41",  x"a4",  x"e8", -- 22D0
         x"9a",  x"dd",  x"be",  x"02",  x"35",  x"28",  x"17",  x"70", -- 22D8
         x"03",  x"8b",  x"07",  x"0f",  x"3e",  x"2a",  x"e8",  x"d1", -- 22E0
         x"e8",  x"f1",  x"19",  x"eb",  x"bd",  x"8e",  x"c0",  x"05", -- 22E8
         x"da",  x"29",  x"7b",  x"3d",  x"46",  x"6e",  x"cd",  x"dd", -- 22F0
         x"2b",  x"13",  x"3e",  x"14",  x"30",  x"a2",  x"41",  x"18", -- 22F8
         x"af",  x"b5",  x"f3",  x"09",  x"4f",  x"00",  x"3f",  x"10", -- 2300
         x"16",  x"ad",  x"f8",  x"28",  x"18",  x"d2",  x"10",  x"2a", -- 2308
         x"08",  x"ba",  x"33",  x"57",  x"09",  x"e5",  x"c3",  x"bc", -- 2310
         x"c7",  x"00",  x"eb",  x"2b",  x"e5",  x"9b",  x"35",  x"b8", -- 2318
         x"b3",  x"d0",  x"c3",  x"88",  x"03",  x"3e",  x"80",  x"d5", -- 2320
         x"4f",  x"3b",  x"c0",  x"c6",  x"22",  x"41",  x"32",  x"c1", -- 2328
         x"83",  x"c9",  x"f0",  x"ab",  x"ca",  x"63",  x"33",  x"00", -- 2330
         x"c3",  x"79",  x"32",  x"04",  x"05",  x"ca",  x"87",  x"33", -- 2338
         x"03",  x"77",  x"2b",  x"04",  x"c3",  x"b2",  x"32",  x"09", -- 2340
         x"cd",  x"03",  x"fa",  x"9a",  x"14",  x"b0",  x"4c",  x"14", -- 2348
         x"c2",  x"04",  x"d1",  x"7b",  x"00",  x"95",  x"3d",  x"12", -- 2350
         x"c1",  x"eb",  x"2a",  x"2b",  x"3d",  x"74",  x"2b",  x"f8", -- 2358
         x"20",  x"7a",  x"cc",  x"85",  x"fe",  x"51",  x"09",  x"04", -- 2360
         x"eb",  x"c9",  x"59",  x"31",  x"24",  x"cd",  x"df",  x"ed", -- 2368
         x"31",  x"05",  x"f5",  x"ed",  x"00",  x"af",  x"3d",  x"cd", -- 2370
         x"87",  x"0d",  x"d2",  x"00",  x"d0",  x"33",  x"23",  x"36", -- 2378
         x"0d",  x"2b",  x"eb",  x"e1",  x"3c",  x"f1",  x"c9",  x"02", -- 2380
         x"97",  x"7c",  x"dd",  x"01",  x"23",  x"31",  x"fe",  x"26", -- 2388
         x"ca",  x"d5",  x"33",  x"da",  x"e7",  x"ca",  x"80",  x"09", -- 2390
         x"21",  x"d0",  x"fe",  x"0d",  x"c8",  x"f5",  x"06",  x"cd", -- 2398
         x"08",  x"0c",  x"ca",  x"f5",  x"37",  x"0f",  x"df",  x"3d", -- 23A0
         x"c1",  x"d8",  x"33",  x"c3",  x"16",  x"21",  x"ff",  x"69", -- 23A8
         x"00",  x"6c",  x"0d",  x"3f",  x"53",  x"74",  x"61",  x"63", -- 23B0
         x"6b",  x"00",  x"20",  x"6f",  x"76",  x"65",  x"72",  x"66", -- 23B8
         x"6c",  x"6f",  x"78",  x"77",  x"a0",  x"74",  x"00",  x"72", -- 23C0
         x"79",  x"20",  x"6d",  x"6f",  x"72",  x"65",  x"20",  x"00", -- 23C8
         x"50",  x"20",  x"73",  x"77",  x"69",  x"74",  x"63",  x"68", -- 23D0
         x"28",  x"65",  x"73",  x"e2",  x"00",  x"cd",  x"a9",  x"28", -- 23D8
         x"3a",  x"f6",  x"3d",  x"a8",  x"f7",  x"31",  x"34",  x"34", -- 23E0
         x"ec",  x"00",  x"00",  x"eb",  x"22",  x"e2",  x"3f",  x"cd", -- 23E8
         x"e3",  x"2f",  x"ad",  x"c7",  x"07",  x"01",  x"48",  x"34", -- 23F0
         x"c5",  x"d5",  x"ec",  x"00",  x"c3",  x"56",  x"04",  x"c1", -- 23F8
         x"01",  x"63",  x"43",  x"0a",  x"cd",  x"4f",  x"0b",  x"72", -- 2400
         x"67",  x"cc",  x"04",  x"cd",  x"2d",  x"9c",  x"2c",  x"69", -- 2408
         x"29",  x"2d",  x"3d",  x"c8",  x"96",  x"20",  x"3a",  x"60", -- 2410
         x"13",  x"7d",  x"c2",  x"5e",  x"34",  x"c9",  x"af",  x"a1", -- 2418
         x"0a",  x"cd",  x"83",  x"3a",  x"47",  x"34",  x"21",  x"cc", -- 2420
         x"f1",  x"cc",  x"d5",  x"af",  x"58",  x"40",  x"aa",  x"b5", -- 2428
         x"2a",  x"47",  x"e5",  x"8d",  x"0d",  x"21",  x"8b",  x"34", -- 2430
         x"dc",  x"b0",  x"b5",  x"36",  x"de",  x"34",  x"d8",  x"61", -- 2438
         x"d1",  x"ce",  x"80",  x"2e",  x"ba",  x"34",  x"3a",  x"eb", -- 2440
         x"3f",  x"b7",  x"c2",  x"3e",  x"a3",  x"34",  x"ec",  x"a3", -- 2448
         x"0b",  x"2a",  x"dd",  x"25",  x"1b",  x"cd",  x"79",  x"39", -- 2450
         x"d0",  x"06",  x"6f",  x"30",  x"af",  x"32",  x"17",  x"d1", -- 2458
         x"d9",  x"3b",  x"e4",  x"10",  x"eb",  x"e9",  x"98",  x"c9", -- 2460
         x"57",  x"3a",  x"b7",  x"2c",  x"ca",  x"ed",  x"66",  x"cd", -- 2468
         x"6d",  x"ca",  x"5a",  x"bd",  x"33",  x"67",  x"51",  x"c5", -- 2470
         x"47",  x"2a",  x"e6",  x"95",  x"1d",  x"2a",  x"e8",  x"03", -- 2478
         x"b7",  x"25",  x"e9",  x"6c",  x"22",  x"05",  x"ff",  x"03", -- 2480
         x"0d",  x"03",  x"15",  x"83",  x"32",  x"0b",  x"62",  x"6b", -- 2488
         x"c3",  x"90",  x"5b",  x"6c",  x"df",  x"5b",  x"ca",  x"bf", -- 2490
         x"6a",  x"4a",  x"83",  x"6e",  x"11",  x"10",  x"35",  x"d5", -- 2498
         x"33",  x"c0",  x"57",  x"ea",  x"3f",  x"c3",  x"3a",  x"0b", -- 24A0
         x"c3",  x"2c",  x"bb",  x"04",  x"78",  x"ca",  x"6f",  x"60", -- 24A8
         x"35",  x"ce",  x"de",  x"44",  x"01",  x"86",  x"ce",  x"b4", -- 24B0
         x"20",  x"c0",  x"b7",  x"f0",  x"4f",  x"e6",  x"00",  x"08", -- 24B8
         x"c2",  x"43",  x"35",  x"79",  x"e6",  x"10",  x"c2",  x"50", -- 24C0
         x"4b",  x"05",  x"20",  x"c2",  x"53",  x"a0",  x"05",  x"40", -- 24C8
         x"c2",  x"60",  x"35",  x"35",  x"c9",  x"3a",  x"3b",  x"3d", -- 24D0
         x"5a",  x"3f",  x"07",  x"3c",  x"60",  x"07",  x"b7",  x"c0", -- 24D8
         x"3a",  x"d8",  x"6a",  x"3c",  x"ee",  x"c3",  x"24",  x"cf", -- 24E0
         x"28",  x"0c",  x"dc",  x"a1",  x"fe",  x"08",  x"a3",  x"eb", -- 24E8
         x"13",  x"c3",  x"35",  x"29",  x"86",  x"fe",  x"ed",  x"05", -- 24F0
         x"b7",  x"f5",  x"09",  x"c2",  x"22",  x"ec",  x"88",  x"c8", -- 24F8
         x"4e",  x"32",  x"4f",  x"94",  x"db",  x"45",  x"95",  x"35", -- 2500
         x"2a",  x"61",  x"0e",  x"e4",  x"90",  x"c4",  x"79",  x"36", -- 2508
         x"00",  x"7e",  x"2b",  x"ac",  x"c4",  x"01",  x"97",  x"04", -- 2510
         x"f1",  x"f5",  x"ca",  x"d1",  x"35",  x"96",  x"cd",  x"86", -- 2518
         x"0b",  x"3c",  x"0c",  x"0e",  x"77",  x"e5",  x"f5",  x"0e", -- 2520
         x"18",  x"f3",  x"2c",  x"7d",  x"2c",  x"36",  x"1b",  x"61", -- 2528
         x"47",  x"c5",  x"8c",  x"1c",  x"71",  x"32",  x"0c",  x"f8", -- 2530
         x"00",  x"ca",  x"29",  x"36",  x"fe",  x"3e",  x"ca",  x"cc", -- 2538
         x"13",  x"c3",  x"c0",  x"10",  x"1d",  x"0b",  x"20",  x"d6", -- 2540
         x"ff",  x"04",  x"f7",  x"00",  x"02",  x"5c",  x"98",  x"01", -- 2548
         x"1c",  x"d5",  x"79",  x"00",  x"01",  x"c3",  x"01",  x"f6", -- 2550
         x"f0",  x"c3",  x"4f",  x"e6",  x"c3",  x"63",  x"80",  x"02", -- 2558
         x"db",  x"e6",  x"08",  x"fd",  x"c3",  x"a7",  x"f8",  x"00", -- 2560
         x"7f",  x"7f",  x"42",  x"41",  x"53",  x"49",  x"43",  x"00", -- 2568
         x"03",  x"cd",  x"2f",  x"e0",  x"c3",  x"0d",  x"c0",  x"0d", -- 2570
         x"22",  x"52",  x"45",  x"40",  x"0f",  x"8c",  x"c0",  x"db", -- 2578
         x"88",  x"f6",  x"80",  x"00",  x"d3",  x"88",  x"dd",  x"7e", -- 2580
         x"04",  x"f6",  x"60",  x"d3",  x"00",  x"86",  x"dd",  x"77", -- 2588
         x"04",  x"c9",  x"ed",  x"5b",  x"a0",  x"01",  x"b7",  x"2a", -- 2590
         x"9c",  x"b7",  x"19",  x"cb",  x"24",  x"60",  x"01",  x"f5", -- 2598
         x"7d",  x"6c",  x"fe",  x"28",  x"30",  x"30",  x"06",  x"23", -- 25A0
         x"67",  x"f1",  x"a7",  x"c9",  x"00",  x"f1",  x"37",  x"c9", -- 25A8
         x"3a",  x"9e",  x"b7",  x"3d",  x"93",  x"18",  x"d8",  x"3a", -- 25B0
         x"9f",  x"05",  x"92",  x"c9",  x"f5",  x"03",  x"cd",  x"5e", -- 25B8
         x"e0",  x"38",  x"eb",  x"3a",  x"2b",  x"00",  x"83",  x"d5", -- 25C0
         x"5f",  x"3a",  x"9d",  x"b7",  x"82",  x"87",  x"c0",  x"00", -- 25C8
         x"6f",  x"26",  x"00",  x"54",  x"29",  x"29",  x"60",  x"19", -- 25D0
         x"43",  x"cb",  x"b7",  x"5f",  x"19",  x"d1",  x"f0",  x"32", -- 25D8
         x"23",  x"e6",  x"c0",  x"4f",  x"f1",  x"d4",  x"04",  x"07", -- 25E0
         x"00",  x"b1",  x"de",  x"08",  x"0f",  x"00",  x"0a",  x"b1", -- 25E8
         x"05",  x"c9",  x"e5",  x"d5",  x"c5",  x"f5",  x"80",  x"62", -- 25F0
         x"eb",  x"21",  x"a6",  x"b7",  x"87",  x"30",  x"02",  x"00", -- 25F8
         x"2e",  x"aa",  x"d6",  x"40",  x"38",  x"04",  x"fe",  x"80", -- 2600
         x"c0",  x"03",  x"c6",  x"40",  x"2c",  x"2c",  x"4e",  x"2c", -- 2608
         x"58",  x"46",  x"46",  x"29",  x"09",  x"7b",  x"a6",  x"78", -- 2610
         x"56",  x"78",  x"42",  x"2b",  x"57",  x"78",  x"58",  x"60", -- 2618
         x"00",  x"a2",  x"b7",  x"cb",  x"57",  x"28",  x"0f",  x"4f", -- 2620
         x"06",  x"00",  x"08",  x"d5",  x"7e",  x"2f",  x"12",  x"23", -- 2628
         x"13",  x"10",  x"00",  x"f9",  x"79",  x"0f",  x"18",  x"14", -- 2630
         x"0f",  x"38",  x"12",  x"11",  x"d5",  x"ed",  x"a0",  x"ad", -- 2638
         x"01",  x"d1",  x"14",  x"1f",  x"80",  x"cf",  x"01",  x"67", -- 2640
         x"ee",  x"00",  x"02",  x"f3",  x"d3",  x"84",  x"3a",  x"a3", -- 2648
         x"b7",  x"12",  x"46",  x"13",  x"30",  x"01",  x"7c",  x"14", -- 2650
         x"fb",  x"f1",  x"c1",  x"d1",  x"48",  x"e1",  x"85",  x"01", -- 2658
         x"08",  x"f5",  x"79",  x"08",  x"41",  x"d2",  x"c7",  x"0a", -- 2660
         x"8c",  x"44",  x"ea",  x"36",  x"e1",  x"22",  x"24",  x"14", -- 2668
         x"00",  x"08",  x"4f",  x"08",  x"3d",  x"20",  x"e1",  x"08", -- 2670
         x"f1",  x"16",  x"08",  x"18",  x"cc",  x"97",  x"2a",  x"21", -- 2678
         x"84",  x"00",  x"66",  x"28",  x"22",  x"cb",  x"00",  x"a6", -- 2680
         x"fe",  x"30",  x"d8",  x"fe",  x"3a",  x"30",  x"04",  x"00", -- 2688
         x"d6",  x"30",  x"18",  x"0a",  x"fe",  x"41",  x"d8",  x"cb", -- 2690
         x"00",  x"af",  x"fe",  x"5b",  x"d0",  x"d6",  x"37",  x"21", -- 2698
         x"df",  x"00",  x"b7",  x"be",  x"d0",  x"87",  x"2a",  x"dd", -- 26A0
         x"b7",  x"18",  x"0c",  x"0c",  x"fe",  x"20",  x"30",  x"c0", -- 26A8
         x"46",  x"5e",  x"20",  x"15",  x"0d",  x"b2",  x"60",  x"b7", -- 26B0
         x"b2",  x"00",  x"00",  x"09",  x"7e",  x"23",  x"66",  x"6f", -- 26B8
         x"e9",  x"7b",  x"e6",  x"00",  x"f8",  x"c6",  x"08",  x"5f", -- 26C0
         x"18",  x"09",  x"cd",  x"6a",  x"01",  x"e0",  x"d8",  x"77", -- 26C8
         x"cd",  x"a3",  x"e0",  x"1c",  x"62",  x"cc",  x"bb",  x"0a", -- 26D0
         x"d0",  x"1e",  x"00",  x"14",  x"cf",  x"10",  x"ba",  x"c0", -- 26D8
         x"2a",  x"a4",  x"0c",  x"b7",  x"e9",  x"2a",  x"99",  x"03", -- 26E0
         x"7b",  x"a7",  x"00",  x"28",  x"02",  x"1d",  x"c9",  x"7a", -- 26E8
         x"a7",  x"c8",  x"15",  x"b4",  x"1f",  x"5f",  x"80",  x"09", -- 26F0
         x"c9",  x"21",  x"45",  x"e2",  x"22",  x"f0",  x"1f",  x"06", -- 26F8
         x"60",  x"e2",  x"18",  x"f7",  x"0a",  x"cd",  x"c1",  x"e1", -- 2700
         x"d5",  x"43",  x"6c",  x"7e",  x"27",  x"29",  x"b8",  x"14", -- 2708
         x"1c",  x"09",  x"30",  x"55",  x"08",  x"43",  x"14",  x"07", -- 2710
         x"38",  x"10",  x"13",  x"0c",  x"0b",  x"42",  x"4b",  x"d1", -- 2718
         x"e3",  x"5e",  x"14",  x"50",  x"59",  x"18",  x"c3",  x"01", -- 2720
         x"36",  x"00",  x"3e",  x"20",  x"42",  x"0c",  x"d1",  x"c9", -- 2728
         x"d5",  x"b5",  x"07",  x"22",  x"46",  x"b4",  x"19",  x"78", -- 2730
         x"25",  x"0e",  x"89",  x"37",  x"f1",  x"4e",  x"37",  x"30", -- 2738
         x"e9",  x"1e",  x"80",  x"82",  x"16",  x"00",  x"c8",  x"d1", -- 2740
         x"aa",  x"e2",  x"30",  x"f1",  x"14",  x"f1",  x"78",  x"f7", -- 2748
         x"0a",  x"19",  x"c9",  x"41",  x"55",  x"23",  x"77",  x"2c", -- 2750
         x"02",  x"01",  x"6a",  x"24",  x"10",  x"ec",  x"ce",  x"81", -- 2758
         x"82",  x"d1",  x"cc",  x"81",  x"28",  x"3d",  x"05",  x"d5", -- 2760
         x"f5",  x"11",  x"00",  x"00",  x"64",  x"40",  x"c8",  x"28", -- 2768
         x"03",  x"00",  x"19",  x"e5",  x"c5",  x"ed",  x"b0",  x"d7", -- 2770
         x"1c",  x"3c",  x"f3",  x"f1",  x"a2",  x"af",  x"50",  x"4f", -- 2778
         x"18",  x"42",  x"cd",  x"44",  x"c5",  x"19",  x"2e",  x"08", -- 2780
         x"19",  x"10",  x"ba",  x"1f",  x"1f",  x"38",  x"60",  x"0b", -- 2788
         x"5c",  x"de",  x"e2",  x"cd",  x"29",  x"e1",  x"f3",  x"05", -- 2790
         x"62",  x"17",  x"d4",  x"07",  x"3b",  x"d1",  x"15",  x"62", -- 2798
         x"89",  x"1a",  x"4f",  x"01",  x"47",  x"4f",  x"af",  x"77", -- 27A0
         x"23",  x"10",  x"fc",  x"ea",  x"2e",  x"0d",  x"d5",  x"2c", -- 27A8
         x"00",  x"0f",  x"5f",  x"38",  x"06",  x"af",  x"e5",  x"cd", -- 27B0
         x"4a",  x"02",  x"e2",  x"e1",  x"cb",  x"0b",  x"38",  x"0c", -- 27B8
         x"a8",  x"2f",  x"c4",  x"aa",  x"0d",  x"b0",  x"08",  x"a6", -- 27C0
         x"a2",  x"d8",  x"a2",  x"d7",  x"d1",  x"a7",  x"01",  x"44", -- 27C8
         x"c5",  x"c9",  x"00",  x"01",  x"0f",  x"0a",  x"21",  x"30", -- 27D0
         x"00",  x"d5",  x"5c",  x"00",  x"cd",  x"2e",  x"f9",  x"3e", -- 27D8
         x"1e",  x"cd",  x"e0",  x"f1",  x"00",  x"3e",  x"03",  x"d3", -- 27E0
         x"8c",  x"3e",  x"10",  x"d1",  x"c3",  x"e7",  x"09",  x"16", -- 27E8
         x"d8",  x"30",  x"21",  x"3b",  x"7e",  x"cd",  x"8e",  x"0a", -- 27F0
         x"e0",  x"77",  x"c9",  x"7e",  x"3b",  x"19",  x"08",  x"ee", -- 27F8
         x"20",  x"3a",  x"08",  x"c9",  x"64",  x"c6",  x"e6",  x"90", -- 2800
         x"ff",  x"81",  x"cd",  x"58",  x"e1",  x"ed",  x"53",  x"94", -- 2808
         x"d7",  x"86",  x"8f",  x"fb",  x"00",  x"f5",  x"3e",  x"23", -- 2810
         x"d3",  x"8f",  x"dd",  x"36",  x"0d",  x"03",  x"00",  x"18", -- 2818
         x"5e",  x"f5",  x"db",  x"8f",  x"0d",  x"66",  x"a7",  x"0d", -- 2820
         x"3e",  x"8f",  x"03",  x"f1",  x"00",  x"fb",  x"b7",  x"28", -- 2828
         x"4d",  x"fe",  x"14",  x"38",  x"49",  x"00",  x"fe",  x"78", -- 2830
         x"30",  x"45",  x"fe",  x"65",  x"30",  x"3d",  x"0f",  x"c6", -- 2838
         x"be",  x"38",  x"39",  x"3c",  x"4d",  x"00",  x"0c",  x"1f", -- 2840
         x"ee",  x"01",  x"dd",  x"6e",  x"0e",  x"dd",  x"31",  x"66", -- 2848
         x"0f",  x"ae",  x"d1",  x"ed",  x"7e",  x"83",  x"42",  x"dd", -- 2850
         x"cb",  x"08",  x"7e",  x"20",  x"90",  x"3d",  x"cc",  x"1a", -- 2858
         x"06",  x"cc",  x"69",  x"d6",  x"40",  x"6b",  x"be",  x"0d", -- 2860
         x"20",  x"1d",  x"f5",  x"18",  x"3a",  x"e0",  x"b7",  x"08", -- 2868
         x"0a",  x"38",  x"11",  x"03",  x"f1",  x"dd",  x"34",  x"0a", -- 2870
         x"18",  x"04",  x"23",  x"00",  x"0c",  x"1e",  x"db",  x"89", -- 2878
         x"d3",  x"89",  x"f1",  x"ed",  x"0c",  x"4d",  x"f1",  x"18", -- 2880
         x"08",  x"6d",  x"0a",  x"00",  x"0c",  x"fe",  x"16",  x"28", -- 2888
         x"09",  x"95",  x"14",  x"0d",  x"3c",  x"c6",  x"2c",  x"18", -- 2890
         x"e5",  x"a3",  x"14",  x"80",  x"a3",  x"01",  x"3e",  x"16", -- 2898
         x"18",  x"eb",  x"e6",  x"36",  x"12",  x"46",  x"c8",  x"11", -- 28A0
         x"0d",  x"d4",  x"f6",  x"cd",  x"ca",  x"29",  x"e3",  x"d0", -- 28A8
         x"0d",  x"86",  x"20",  x"08",  x"fe",  x"03",  x"37",  x"6b", -- 28B0
         x"c8",  x"d9",  x"b0",  x"c8",  x"53",  x"57",  x"49",  x"00", -- 28B8
         x"54",  x"43",  x"48",  x"01",  x"53",  x"cd",  x"04",  x"e4", -- 28C0
         x"05",  x"7d",  x"cd",  x"59",  x"f3",  x"7c",  x"00",  x"03", -- 28C8
         x"7a",  x"cd",  x"76",  x"f3",  x"c3",  x"6b",  x"f3",  x"0c", -- 28D0
         x"26",  x"b8",  x"0e",  x"80",  x"aa",  x"1a",  x"02",  x"a0", -- 28D8
         x"00",  x"56",  x"ed",  x"60",  x"c9",  x"72",  x"7d",  x"fe", -- 28E0
         x"00",  x"05",  x"38",  x"14",  x"ed",  x"51",  x"18",  x"f3", -- 28E8
         x"e6",  x"00",  x"f5",  x"cb",  x"42",  x"28",  x"5c",  x"cb", -- 28F0
         x"cf",  x"cb",  x"00",  x"4a",  x"28",  x"56",  x"cb",  x"df", -- 28F8
         x"18",  x"52",  x"fe",  x"14",  x"04",  x"38",  x"18",  x"f9", -- 2900
         x"c5",  x"e6",  x"fc",  x"0a",  x"16",  x"08",  x"cb",  x"c7", -- 2908
         x"16",  x"74",  x"02",  x"1c",  x"83",  x"fb",  x"88",  x"99", -- 2910
         x"18",  x"38",  x"64",  x"38",  x"24",  x"81",  x"a7",  x"e6", -- 2918
         x"9f",  x"22",  x"1a",  x"ef",  x"46",  x"1a",  x"f7",  x"b5", -- 2920
         x"14",  x"fe",  x"20",  x"f6",  x"10",  x"cb",  x"52",  x"20", -- 2928
         x"c1",  x"dc",  x"10",  x"95",  x"80",  x"11",  x"85",  x"18", -- 2930
         x"10",  x"9b",  x"65",  x"38",  x"0f",  x"c3",  x"e5",  x"25", -- 2938
         x"cb",  x"bf",  x"37",  x"21",  x"ff",  x"c9",  x"06",  x"26", -- 2940
         x"ff",  x"c9",  x"fe",  x"01",  x"10",  x"da",  x"28",  x"1b", -- 2948
         x"e4",  x"13",  x"97",  x"28",  x"06",  x"ee",  x"cb",  x"d7", -- 2950
         x"18",  x"ea",  x"aa",  x"00",  x"4a",  x"55",  x"4d",  x"50", -- 2958
         x"01",  x"30",  x"7d",  x"47",  x"95",  x"00",  x"ed",  x"78", -- 2960
         x"3c",  x"ca",  x"61",  x"f3",  x"3e",  x"ff",  x"c0",  x"a1", -- 2968
         x"68",  x"77",  x"18",  x"f3",  x"ed",  x"79",  x"28",  x"e6", -- 2970
         x"7e",  x"c3",  x"15",  x"b4",  x"b7",  x"f3",  x"85",  x"03", -- 2978
         x"40",  x"e6",  x"df",  x"3d",  x"52",  x"fb",  x"84",  x"99", -- 2980
         x"22",  x"cf",  x"ed",  x"06",  x"fd",  x"f1",  x"22",  x"cd", -- 2988
         x"05",  x"d6",  x"59",  x"e1",  x"d1",  x"14",  x"d3",  x"8d", -- 2990
         x"f9",  x"03",  x"8e",  x"18",  x"28",  x"ab",  x"10",  x"02", -- 2998
         x"fe",  x"cd",  x"2b",  x"33",  x"e5",  x"2a",  x"18",  x"22", -- 29A0
         x"b9",  x"a1",  x"8e",  x"24",  x"94",  x"8f",  x"21",  x"80", -- 29A8
         x"02",  x"b7",  x"af",  x"2d",  x"77",  x"20",  x"fc",  x"9b", -- 29B0
         x"46",  x"9f",  x"3c",  x"cd",  x"f8",  x"0b",  x"a3",  x"1c", -- 29B8
         x"03",  x"01",  x"5e",  x"30",  x"28",  x"06",  x"bb",  x"a0", -- 29C0
         x"8d",  x"50",  x"89",  x"0f",  x"4e",  x"20",  x"fa",  x"03", -- 29C8
         x"3e",  x"47",  x"d3",  x"8e",  x"3e",  x"0c",  x"03",  x"58", -- 29D0
         x"c9",  x"67",  x"60",  x"cd",  x"bb",  x"50",  x"e4",  x"4a", -- 29D8
         x"00",  x"01",  x"00",  x"65",  x"10",  x"90",  x"99",  x"ca", -- 29E0
         x"3e",  x"87",  x"98",  x"5f",  x"3e",  x"2f",  x"03",  x"fb", -- 29E8
         x"57",  x"5f",  x"01",  x"cd",  x"80",  x"e5",  x"ed",  x"a1", -- 29F0
         x"ea",  x"3a",  x"9a",  x"f9",  x"7e",  x"89",  x"86",  x"02", -- 29F8
         x"e6",  x"4d",  x"05",  x"6e",  x"05",  x"dc",  x"41",  x"06", -- 2A00
         x"06",  x"80",  x"7e",  x"43",  x"0b",  x"79",  x"86",  x"4f", -- 2A08
         x"a2",  x"45",  x"f6",  x"62",  x"08",  x"e2",  x"83",  x"18", -- 2A10
         x"e5",  x"5d",  x"54",  x"98",  x"65",  x"32",  x"c9",  x"c5", -- 2A18
         x"40",  x"8d",  x"cb",  x"09",  x"1e",  x"d3",  x"cd",  x"38", -- 2A20
         x"18",  x"1e",  x"2f",  x"dc",  x"04",  x"10",  x"f2",  x"c1", -- 2A28
         x"3c",  x"1e",  x"5d",  x"1e",  x"37",  x"72",  x"00",  x"cd", -- 2A30
         x"40",  x"00",  x"a7",  x"78",  x"53",  x"90",  x"af",  x"b4", -- 2A38
         x"e4",  x"3e",  x"19",  x"83",  x"d3",  x"8a",  x"ae",  x"96", -- 2A40
         x"06",  x"16",  x"d9",  x"60",  x"cd",  x"1a",  x"e6",  x"38", -- 2A48
         x"f5",  x"01",  x"fe",  x"ba",  x"cd",  x"ed",  x"e5",  x"38", -- 2A50
         x"ee",  x"86",  x"2d",  x"06",  x"02",  x"af",  x"4f",  x"c4", -- 2A58
         x"38",  x"14",  x"2d",  x"e6",  x"fe",  x"19",  x"5d",  x"30", -- 2A60
         x"f2",  x"0f",  x"cd",  x"39",  x"b7",  x"1d",  x"25",  x"10", -- 2A68
         x"02",  x"71",  x"2d",  x"79",  x"94",  x"0f",  x"15",  x"77", -- 2A70
         x"80",  x"75",  x"98",  x"4d",  x"0d",  x"7d",  x"f0",  x"78", -- 2A78
         x"0f",  x"17",  x"96",  x"0d",  x"c6",  x"67",  x"ff",  x"eb", -- 2A80
         x"83",  x"b8",  x"03",  x"56",  x"50",  x"fb",  x"f9",  x"b3", -- 2A88
         x"ef",  x"e9",  x"df",  x"ff",  x"fc",  x"0e",  x"e9",  x"6c", -- 2A90
         x"c9",  x"2a",  x"76",  x"b6",  x"04",  x"f3",  x"d1",  x"c2", -- 2A98
         x"0e",  x"a2",  x"c2",  x"8e",  x"8a",  x"5b",  x"3e",  x"07", -- 2AA0
         x"fa",  x"07",  x"a3",  x"03",  x"a6",  x"c4",  x"ef",  x"77", -- 2AA8
         x"17",  x"f5",  x"30",  x"2a",  x"24",  x"a1",  x"d1",  x"f6", -- 2AB0
         x"4f",  x"1a",  x"0e",  x"81",  x"6c",  x"c9",  x"b1",  x"08", -- 2AB8
         x"b0",  x"9e",  x"60",  x"03",  x"9e",  x"d8",  x"02",  x"3f", -- 2AC0
         x"cb",  x"1b",  x"15",  x"20",  x"f2",  x"80",  x"0d",  x"7b", -- 2AC8
         x"c9",  x"78",  x"d6",  x"09",  x"38",  x"02",  x"4f",  x"fe", -- 2AD0
         x"1b",  x"30",  x"4b",  x"07",  x"9b",  x"f5",  x"e7",  x"67", -- 2AD8
         x"ba",  x"d1",  x"60",  x"b7",  x"c8",  x"7e",  x"fe",  x"df", -- 2AE0
         x"e2",  x"fe",  x"90",  x"87",  x"e1",  x"ca",  x"62",  x"97", -- 2AE8
         x"ae",  x"fd",  x"60",  x"03",  x"e8",  x"2e",  x"35",  x"3c", -- 2AF0
         x"32",  x"06",  x"e5",  x"28",  x"ea",  x"cd",  x"95",  x"ec", -- 2AF8
         x"0a",  x"e1",  x"32",  x"7e",  x"03",  x"20",  x"00",  x"28", -- 2B00
         x"1d",  x"fe",  x"e2",  x"ca",  x"9b",  x"e6",  x"cd",  x"06", -- 2B08
         x"bd",  x"c8",  x"cd",  x"14",  x"eb",  x"0f",  x"3b",  x"df", -- 2B10
         x"ac",  x"ed",  x"4b",  x"0c",  x"01",  x"30",  x"eb",  x"18", -- 2B18
         x"f1",  x"c3",  x"48",  x"c3",  x"65",  x"0a",  x"fa",  x"ea", -- 2B20
         x"80",  x"17",  x"25",  x"cd",  x"cc",  x"c8",  x"2c",  x"fe", -- 2B28
         x"e0",  x"25",  x"20",  x"ea",  x"2a",  x"a0",  x"0d",  x"3b", -- 2B30
         x"cd",  x"03",  x"cb",  x"25",  x"3a",  x"7e",  x"4f",  x"6c", -- 2B38
         x"91",  x"4f",  x"c1",  x"e7",  x"4a",  x"18",  x"a3",  x"1c", -- 2B40
         x"00",  x"18",  x"e8",  x"79",  x"fe",  x"62",  x"ca",  x"4b", -- 2B48
         x"ea",  x"00",  x"fe",  x"6e",  x"ca",  x"c3",  x"ec",  x"fe", -- 2B50
         x"7c",  x"ca",  x"00",  x"a1",  x"ed",  x"fe",  x"76",  x"ca", -- 2B58
         x"c4",  x"ed",  x"d6",  x"39",  x"3e",  x"38",  x"fe",  x"00", -- 2B60
         x"07",  x"30",  x"ab",  x"eb",  x"01",  x"b2",  x"fd",  x"e1", -- 2B68
         x"1c",  x"6f",  x"09",  x"4e",  x"e9",  x"85",  x"69",  x"e5", -- 2B70
         x"eb",  x"c9",  x"06",  x"46",  x"28",  x"cd",  x"21",  x"d4", -- 2B78
         x"e0",  x"cc",  x"d6",  x"54",  x"3a",  x"cd",  x"06",  x"cd", -- 2B80
         x"db",  x"c8",  x"f1",  x"e5",  x"0b",  x"30",  x"01",  x"d3", -- 2B88
         x"23",  x"23",  x"5e",  x"23",  x"56",  x"c1",  x"b3",  x"f7", -- 2B90
         x"d5",  x"f1",  x"77",  x"b9",  x"a9",  x"2d",  x"b8",  x"f8", -- 2B98
         x"40",  x"79",  x"05",  x"28",  x"05",  x"81",  x"38",  x"1a", -- 2BA0
         x"2b",  x"10",  x"fb",  x"9b",  x"0e",  x"00",  x"c5",  x"cd", -- 2BA8
         x"94",  x"1a",  x"c1",  x"1c",  x"cd",  x"98",  x"c9",  x"e3", -- 2BB0
         x"7c",  x"c7",  x"02",  x"6f",  x"24",  x"25",  x"d2",  x"00", -- 2BB8
         x"28",  x"07",  x"cd",  x"f2",  x"d2",  x"e4",  x"ef",  x"18", -- 2BC0
         x"f4",  x"c0",  x"03",  x"d1",  x"cd",  x"02",  x"d3",  x"c3", -- 2BC8
         x"a9",  x"03",  x"d1",  x"1e",  x"1c",  x"c3",  x"56",  x"c3", -- 2BD0
         x"9b",  x"0d",  x"b7",  x"80",  x"22",  x"54",  x"03",  x"2a", -- 2BD8
         x"5f",  x"03",  x"3b",  x"f5",  x"e5",  x"53",  x"dd",  x"a0", -- 2BE0
         x"22",  x"4e",  x"03",  x"22",  x"3b",  x"52",  x"03",  x"a4", -- 2BE8
         x"02",  x"d7",  x"03",  x"1b",  x"1b",  x"e1",  x"e5",  x"c0", -- 2BF0
         x"11",  x"cd",  x"89",  x"c6",  x"e3",  x"20",  x"f4",  x"4c", -- 2BF8
         x"d1",  x"1e",  x"50",  x"1c",  x"03",  x"06",  x"04",  x"96", -- 2C00
         x"67",  x"24",  x"e3",  x"28",  x"86",  x"5b",  x"c6",  x"03", -- 2C08
         x"f5",  x"7a",  x"b3",  x"ca",  x"67",  x"cf",  x"d0",  x"e3", -- 2C10
         x"73",  x"23",  x"72",  x"78",  x"23",  x"d4",  x"f5",  x"7d", -- 2C18
         x"05",  x"66",  x"0b",  x"03",  x"aa",  x"18",  x"9a",  x"90", -- 2C20
         x"c2",  x"69",  x"ea",  x"2a",  x"fe",  x"2b",  x"47",  x"29", -- 2C28
         x"9f",  x"3f",  x"da",  x"23",  x"62",  x"9e",  x"08",  x"be", -- 2C30
         x"c4",  x"9a",  x"9d",  x"28",  x"cf",  x"f8",  x"1e",  x"e1", -- 2C38
         x"c5",  x"17",  x"1b",  x"21",  x"ca",  x"b6",  x"8c",  x"4d", -- 2C40
         x"60",  x"69",  x"e9",  x"00",  x"46",  x"78",  x"b1",  x"28", -- 2C48
         x"b8",  x"23",  x"9a",  x"6b",  x"94",  x"35",  x"23",  x"17", -- 2C50
         x"20",  x"65",  x"e6",  x"70",  x"29",  x"23",  x"80",  x"87", -- 2C58
         x"19",  x"38",  x"c0",  x"0c",  x"cd",  x"27",  x"c3",  x"22", -- 2C60
         x"08",  x"af",  x"2b",  x"78",  x"77",  x"01",  x"95",  x"2d", -- 2C68
         x"eb",  x"6c",  x"3d",  x"ce",  x"e8",  x"01",  x"eb",  x"61", -- 2C70
         x"2a",  x"a9",  x"40",  x"af",  x"e1",  x"a1",  x"41",  x"23", -- 2C78
         x"c5",  x"01",  x"8d",  x"08",  x"7e",  x"12",  x"0a",  x"14", -- 2C80
         x"13",  x"21",  x"06",  x"13",  x"2a",  x"98",  x"0e",  x"ed", -- 2C88
         x"4b",  x"d9",  x"2a",  x"09",  x"1f",  x"85",  x"51",  x"2b", -- 2C90
         x"7c",  x"b5",  x"8a",  x"53",  x"d5",  x"12",  x"e1",  x"87", -- 2C98
         x"04",  x"e5",  x"b8",  x"30",  x"6f",  x"a6",  x"3c",  x"28", -- 2CA0
         x"79",  x"26",  x"76",  x"b4",  x"80",  x"ef",  x"fe",  x"88", -- 2CA8
         x"28",  x"2a",  x"fe",  x"8c",  x"cd",  x"0c",  x"fe",  x"8b", -- 2CB0
         x"a4",  x"c7",  x"fe",  x"d4",  x"28",  x"c3",  x"c0",  x"a9", -- 2CB8
         x"20",  x"e7",  x"cd",  x"87",  x"00",  x"c9",  x"7b",  x"b2", -- 2CC0
         x"c4",  x"ae",  x"e8",  x"c4",  x"e0",  x"0a",  x"e8",  x"18", -- 2CC8
         x"db",  x"2b",  x"7e",  x"b0",  x"7d",  x"e1",  x"e1",  x"c3", -- 2CD0
         x"8a",  x"48",  x"c4",  x"19",  x"28",  x"24",  x"c7",  x"cd", -- 2CD8
         x"1b",  x"c8",  x"fa",  x"2c",  x"20",  x"1a",  x"bc",  x"18", -- 2CE0
         x"ec",  x"98",  x"8d",  x"11",  x"ff",  x"ff",  x"91",  x"85", -- 2CE8
         x"c4",  x"d1",  x"03",  x"61",  x"00",  x"d3",  x"e1",  x"7a", -- 2CF0
         x"99",  x"80",  x"5f",  x"e5",  x"b6",  x"28",  x"16",  x"7e", -- 2CF8
         x"2b",  x"6e",  x"50",  x"67",  x"d5",  x"0a",  x"28",  x"0a", -- 2D00
         x"2a",  x"8c",  x"00",  x"44",  x"4d",  x"e1",  x"23",  x"37", -- 2D08
         x"18",  x"e7",  x"b5",  x"79",  x"b7",  x"47",  x"8c",  x"e1", -- 2D10
         x"bd",  x"80",  x"53",  x"ed",  x"52",  x"e5",  x"c1",  x"62", -- 2D18
         x"6b",  x"1b",  x"65",  x"1a",  x"44",  x"28",  x"0b",  x"71", -- 2D20
         x"88",  x"07",  x"c5",  x"f1",  x"c0",  x"b0",  x"d1",  x"99", -- 2D28
         x"4d",  x"eb",  x"d1",  x"b1",  x"0c",  x"af",  x"06",  x"98", -- 2D30
         x"61",  x"d6",  x"cd",  x"3a",  x"34",  x"d8",  x"d3",  x"c2", -- 2D38
         x"d3",  x"80",  x"a4",  x"0f",  x"c5",  x"cc",  x"8e",  x"09", -- 2D40
         x"54",  x"0e",  x"5d",  x"2b",  x"ed",  x"b8",  x"ea",  x"83", -- 2D48
         x"a0",  x"c1",  x"18",  x"ed",  x"29",  x"50",  x"5b",  x"d2", -- 2D50
         x"94",  x"93",  x"c4",  x"b7",  x"2d",  x"b6",  x"a1",  x"ac", -- 2D58
         x"94",  x"4e",  x"13",  x"13",  x"83",  x"f7",  x"52",  x"e1", -- 2D60
         x"23",  x"83",  x"2d",  x"23",  x"20",  x"fb",  x"c1",  x"e3", -- 2D68
         x"61",  x"28",  x"c9",  x"c8",  x"a3",  x"85",  x"ca",  x"42", -- 2D70
         x"c4",  x"12",  x"92",  x"d5",  x"82",  x"09",  x"e1",  x"c0", -- 2D78
         x"eb",  x"e5",  x"80",  x"a3",  x"d2",  x"4d",  x"c1",  x"a6", -- 2D80
         x"f5",  x"9a",  x"9e",  x"be",  x"c6",  x"08",  x"c1",  x"c3", -- 2D88
         x"50",  x"1d",  x"be",  x"15",  x"c8",  x"20",  x"0f",  x"90", -- 2D90
         x"47",  x"30",  x"fb",  x"ac",  x"23",  x"c8",  x"fe",  x"0a", -- 2D98
         x"eb",  x"26",  x"c3",  x"d8",  x"f4",  x"f3",  x"6f",  x"4f", -- 2DA0
         x"82",  x"1e",  x"1e",  x"d5",  x"9e",  x"15",  x"f0",  x"29", -- 2DA8
         x"1a",  x"c1",  x"25",  x"30",  x"0a",  x"1b",  x"57",  x"03", -- 2DB0
         x"1b",  x"8c",  x"61",  x"e5",  x"c9",  x"06",  x"01",  x"58", -- 2DB8
         x"35",  x"a8",  x"d3",  x"26",  x"47",  x"9a",  x"6a",  x"80", -- 2DC0
         x"dc",  x"26",  x"10",  x"f7",  x"5b",  x"c9",  x"12",  x"65", -- 2DC8
         x"61",  x"c2",  x"13",  x"e3",  x"21",  x"f6",  x"b9",  x"91", -- 2DD0
         x"f2",  x"23",  x"67",  x"8b",  x"71",  x"0e",  x"d3",  x"0b", -- 2DD8
         x"80",  x"0a",  x"57",  x"cd",  x"18",  x"f0",  x"fe",  x"28", -- 2DE0
         x"30",  x"05",  x"4d",  x"3a",  x"f8",  x"b9",  x"5f",  x"03", -- 2DE8
         x"07",  x"45",  x"7a",  x"93",  x"38",  x"41",  x"81",  x"6f", -- 2DF0
         x"c7",  x"40",  x"7b",  x"32",  x"9c",  x"b7",  x"3a",  x"f7", -- 2DF8
         x"57",  x"b9",  x"fc",  x"85",  x"32",  x"57",  x"3a",  x"f6", -- 2E00
         x"e5",  x"07",  x"b5",  x"4d",  x"1b",  x"25",  x"1b",  x"9f", -- 2E08
         x"47",  x"1b",  x"9d",  x"b7",  x"ad",  x"5f",  x"64",  x"39", -- 2E10
         x"99",  x"bf",  x"01",  x"22",  x"fc",  x"27",  x"b1",  x"1e", -- 2E18
         x"76",  x"22",  x"31",  x"cb",  x"7e",  x"fe",  x"0c",  x"cd", -- 2E20
         x"1b",  x"f0",  x"d7",  x"68",  x"04",  x"18",  x"2c",  x"d1", -- 2E28
         x"d7",  x"81",  x"cd",  x"d1",  x"a8",  x"f4",  x"1e",  x"10", -- 2E30
         x"c3",  x"c3",  x"9a",  x"8f",  x"50",  x"cd",  x"e3",  x"11", -- 2E38
         x"f3",  x"62",  x"cd",  x"82",  x"6f",  x"f7",  x"ac",  x"29", -- 2E40
         x"66",  x"80",  x"d0",  x"03",  x"05",  x"3e",  x"bf",  x"bc", -- 2E48
         x"38",  x"07",  x"b0",  x"e4",  x"c3",  x"e9",  x"d3",  x"b6", -- 2E50
         x"c5",  x"7f",  x"6c",  x"d6",  x"30",  x"93",  x"2f",  x"11", -- 2E58
         x"1f",  x"99",  x"0b",  x"20",  x"2f",  x"dd",  x"7a",  x"41", -- 2E60
         x"50",  x"d9",  x"15",  x"0f",  x"00",  x"e6",  x"60",  x"b8", -- 2E68
         x"b7",  x"9f",  x"c3",  x"53",  x"53",  x"f9",  x"a7",  x"9d", -- 2E70
         x"cb",  x"4f",  x"dd",  x"d3",  x"a7",  x"89",  x"20",  x"c6", -- 2E78
         x"d5",  x"03",  x"86",  x"83",  x"06",  x"22",  x"a3",  x"01", -- 2E80
         x"11",  x"ec",  x"b9",  x"01",  x"be",  x"d7",  x"bc",  x"56", -- 2E88
         x"88",  x"16",  x"94",  x"0c",  x"20",  x"94",  x"2c",  x"8e", -- 2E90
         x"32",  x"78",  x"42",  x"eb",  x"9a",  x"b4",  x"de",  x"8c", -- 2E98
         x"9d",  x"cb",  x"38",  x"be",  x"cb",  x"e4",  x"21",  x"19", -- 2EA0
         x"cd",  x"d3",  x"e6",  x"26",  x"37",  x"31",  x"11",  x"e4", -- 2EA8
         x"29",  x"34",  x"bd",  x"28",  x"b1",  x"bf",  x"68",  x"59", -- 2EB0
         x"b8",  x"db",  x"8d",  x"0e",  x"70",  x"80",  x"f2",  x"f6", -- 2EB8
         x"cb",  x"5a",  x"27",  x"01",  x"57",  x"78",  x"8e",  x"0b", -- 2EC0
         x"e6",  x"07",  x"18",  x"12",  x"19",  x"11",  x"08",  x"30", -- 2EC8
         x"dc",  x"24",  x"13",  x"f8",  x"b2",  x"ef",  x"dd",  x"20", -- 2ED0
         x"fc",  x"aa",  x"c2",  x"8b",  x"29",  x"07",  x"c8",  x"6c", -- 2ED8
         x"82",  x"d3",  x"f7",  x"11",  x"eb",  x"99",  x"be",  x"e9", -- 2EE0
         x"30",  x"9f",  x"20",  x"30",  x"3d",  x"ba",  x"38",  x"48", -- 2EE8
         x"9e",  x"8c",  x"79",  x"13",  x"d1",  x"4f",  x"a5",  x"14", -- 2EF0
         x"9e",  x"14",  x"0d",  x"b9",  x"38",  x"89",  x"79",  x"0c", -- 2EF8
         x"a0",  x"64",  x"47",  x"7a",  x"23",  x"8b",  x"4c",  x"e5", -- 2F00
         x"8e",  x"33",  x"0f",  x"3e",  x"e4",  x"26",  x"7b",  x"ad", -- 2F08
         x"f9",  x"f0",  x"05",  x"2a",  x"c2",  x"03",  x"77",  x"3a", -- 2F10
         x"b1",  x"af",  x"b6",  x"0d",  x"bc",  x"ac",  x"3a",  x"2b", -- 2F18
         x"82",  x"b7",  x"de",  x"85",  x"42",  x"d4",  x"d8",  x"f1", -- 2F20
         x"0b",  x"c5",  x"94",  x"b9",  x"73",  x"ef",  x"d2",  x"93", -- 2F28
         x"c1",  x"83",  x"1c",  x"18",  x"f3",  x"5f",  x"10",  x"20", -- 2F30
         x"14",  x"f8",  x"42",  x"1e",  x"35",  x"c1",  x"8b",  x"8f", -- 2F38
         x"bc",  x"3d",  x"33",  x"6c",  x"88",  x"63",  x"7b",  x"21", -- 2F40
         x"d3",  x"89",  x"72",  x"ce",  x"92",  x"40",  x"7e",  x"cd", -- 2F48
         x"10",  x"ec",  x"1e",  x"32",  x"30",  x"c1",  x"5a",  x"01", -- 2F50
         x"1d",  x"8d",  x"d7",  x"da",  x"be",  x"c8",  x"ed",  x"7d", -- 2F58
         x"87",  x"a6",  x"cd",  x"d7",  x"09",  x"06",  x"7e",  x"d6", -- 2F60
         x"b7",  x"17",  x"00",  x"c3",  x"62",  x"78",  x"da",  x"36", -- 2F68
         x"f5",  x"16",  x"12",  x"e5",  x"48",  x"90",  x"28",  x"38", -- 2F70
         x"47",  x"92",  x"93",  x"44",  x"e1",  x"d5",  x"c5",  x"b3", -- 2F78
         x"a7",  x"ab",  x"b5",  x"e5",  x"0a",  x"b7",  x"18",  x"1f", -- 2F80
         x"17",  x"72",  x"cb",  x"c1",  x"7a",  x"4f",  x"10",  x"dd", -- 2F88
         x"83",  x"1a",  x"be",  x"28",  x"12",  x"23",  x"bf",  x"41", -- 2F90
         x"f9",  x"af",  x"e1",  x"d9",  x"00",  x"91",  x"87",  x"c3", -- 2F98
         x"c0",  x"d0",  x"c3",  x"9b",  x"1b",  x"a8",  x"31",  x"2b", -- 2FA0
         x"14",  x"28",  x"0e",  x"13",  x"a9",  x"71",  x"11",  x"20", -- 2FA8
         x"f4",  x"44",  x"8b",  x"0d",  x"c7",  x"be",  x"0d",  x"07", -- 2FB0
         x"e1",  x"20",  x"d8",  x"18",  x"01",  x"0c",  x"b6",  x"00", -- 2FB8
         x"a7",  x"a6",  x"06",  x"7d",  x"18",  x"d0",  x"1e",  x"28", -- 2FC0
         x"f7",  x"61",  x"1e",  x"29",  x"18",  x"0c",  x"40",  x"81", -- 2FC8
         x"a7",  x"fc",  x"f7",  x"fe",  x"0d",  x"0a",  x"30",  x"52", -- 2FD0
         x"1e",  x"39",  x"cc",  x"00",  x"1e",  x"3a",  x"18",  x"f9", -- 2FD8
         x"9e",  x"a1",  x"a8",  x"e9",  x"7a",  x"9f",  x"06",  x"6f", -- 2FE0
         x"3e",  x"02",  x"1e",  x"26",  x"b8",  x"16",  x"8a",  x"91", -- 2FE8
         x"47",  x"f7",  x"16",  x"ec",  x"1e",  x"e4",  x"d6",  x"1e", -- 2FF0
         x"d3",  x"1d",  x"b8",  x"24",  x"23",  x"0d",  x"59",  x"30", -- 2FF8
         x"0d",  x"01",  x"78",  x"32",  x"8b",  x"75",  x"bf",  x"9b", -- 3000
         x"a9",  x"49",  x"cc",  x"a0",  x"0c",  x"fe",  x"4f",  x"20", -- 3008
         x"1e",  x"f1",  x"c5",  x"23",  x"0b",  x"ca",  x"cf",  x"ea", -- 3010
         x"25",  x"58",  x"18",  x"e6",  x"03",  x"c1",  x"e8",  x"06", -- 3018
         x"17",  x"81",  x"f5",  x"3d",  x"37",  x"37",  x"1b",  x"cb", -- 3020
         x"10",  x"3d",  x"df",  x"1b",  x"21",  x"07",  x"e1",  x"80", -- 3028
         x"a8",  x"77",  x"f1",  x"e1",  x"cb",  x"f7",  x"d5",  x"37", -- 3030
         x"5f",  x"16",  x"88",  x"00",  x"0e",  x"e0",  x"d1",  x"c9", -- 3038
         x"ed",  x"5f",  x"32",  x"1d",  x"37",  x"03",  x"c9",  x"8f", -- 3040
         x"a5",  x"3f",  x"19",  x"00",  x"3e",  x"c6",  x"cd",  x"25", -- 3048
         x"de",  x"cd",  x"c8",  x"dd",  x"30",  x"c8",  x"3e",  x"80", -- 3050
         x"0e",  x"b2",  x"dc",  x"21",  x"ea",  x"bf",  x"70",  x"89", -- 3058
         x"50",  x"dd",  x"94",  x"03",  x"5f",  x"de",  x"3a",  x"09", -- 3060
         x"03",  x"4e",  x"88",  x"16",  x"a2",  x"e0",  x"c0",  x"15", -- 3068
         x"01",  x"3e",  x"04",  x"18",  x"03",  x"01",  x"2c",  x"3f", -- 3070
         x"03",  x"98",  x"bb",  x"ba",  x"b2",  x"e0",  x"59",  x"7b", -- 3078
         x"c0",  x"2f",  x"7a",  x"04",  x"96",  x"12",  x"0c",  x"e3", -- 3080
         x"ca",  x"e4",  x"f2",  x"1a",  x"e4",  x"59",  x"e7",  x"9e", -- 3088
         x"22",  x"d1",  x"d5",  x"d5",  x"24",  x"90",  x"91",  x"a7", -- 3090
         x"3e",  x"00",  x"0b",  x"20",  x"06",  x"21",  x"9d",  x"ce", -- 3098
         x"31",  x"47",  x"21",  x"a1",  x"6b",  x"06",  x"80",  x"ce", -- 30A0
         x"04",  x"e3",  x"a7",  x"c1",  x"a7",  x"ec",  x"ab",  x"14", -- 30A8
         x"dd",  x"62",  x"6a",  x"e0",  x"7e",  x"90",  x"e9",  x"c3", -- 30B0
         x"8b",  x"00",  x"eb",  x"9a",  x"e1",  x"6e",  x"f9",  x"7f", -- 30B8
         x"f9",  x"8c",  x"00",  x"f9",  x"9b",  x"f9",  x"8d",  x"f8", -- 30C0
         x"9f",  x"f8",  x"aa",  x"00",  x"f9",  x"0f",  x"e3",  x"b2", -- 30C8
         x"f9",  x"b9",  x"f9",  x"00",  x"06",  x"03",  x"c0",  x"20", -- 30D0
         x"99",  x"c1",  x"bf",  x"a3",  x"4c",  x"58",  x"33",  x"04", -- 30D8
         x"13",  x"00",  x"42",  x"00",  x"2f",  x"00",  x"30",  x"00", -- 30E0
         x"05",  x"09",  x"00",  x"77",  x"33",  x"66",  x"00",  x"0f", -- 30E8
         x"36",  x"36",  x"fe",  x"6c",  x"fe",  x"d8",  x"66",  x"d8", -- 30F0
         x"91",  x"3e",  x"3b",  x"6c",  x"3e",  x"8c",  x"00",  x"7e", -- 30F8
         x"18",  x"00",  x"c6",  x"cc",  x"18",  x"30",  x"66",  x"00", -- 3100
         x"c6",  x"00",  x"38",  x"6c",  x"38",  x"76",  x"dc",  x"cc", -- 3108
         x"0e",  x"76",  x"00",  x"1c",  x"0c",  x"12",  x"f6",  x"00", -- 3110
         x"14",  x"60",  x"00",  x"30",  x"eb",  x"0b",  x"03",  x"00", -- 3118
         x"f0",  x"0b",  x"10",  x"66",  x"3c",  x"ff",  x"3c",  x"bd", -- 3120
         x"42",  x"4d",  x"fc",  x"cd",  x"02",  x"5c",  x"29",  x"2c", -- 3128
         x"fe",  x"00",  x"12",  x"6c",  x"00",  x"78",  x"06",  x"12", -- 3130
         x"2d",  x"c0",  x"80",  x"00",  x"01",  x"7c",  x"c6",  x"ce", -- 3138
         x"de",  x"f6",  x"e6",  x"7c",  x"ab",  x"12",  x"70",  x"7f", -- 3140
         x"32",  x"01",  x"00",  x"78",  x"cc",  x"0c",  x"38",  x"60", -- 3148
         x"cc",  x"b0",  x"07",  x"fc",  x"1e",  x"78",  x"0c",  x"cc", -- 3150
         x"78",  x"c0",  x"3a",  x"3c",  x"6c",  x"cc",  x"fe",  x"0c", -- 3158
         x"1e",  x"c5",  x"0f",  x"c0",  x"f8",  x"0c",  x"fb",  x"0f", -- 3160
         x"1c",  x"08",  x"cc",  x"07",  x"ff",  x"0f",  x"27",  x"21", -- 3168
         x"00",  x"fb",  x"2f",  x"0c",  x"02",  x"b6",  x"07",  x"7c", -- 3170
         x"11",  x"70",  x"97",  x"5c",  x"02",  x"9d",  x"07",  x"60", -- 3178
         x"76",  x"65",  x"9f",  x"1d",  x"00",  x"55",  x"53",  x"05", -- 3180
         x"5d",  x"0b",  x"79",  x"fd",  x"67",  x"06",  x"20",  x"37", -- 3188
         x"7f",  x"de",  x"00",  x"c0",  x"3f",  x"fb",  x"6d",  x"40", -- 3190
         x"53",  x"cc",  x"23",  x"1f",  x"66",  x"66",  x"7c",  x"02", -- 3198
         x"29",  x"83",  x"c3",  x"c0",  x"00",  x"c0",  x"cb",  x"00", -- 31A0
         x"f8",  x"63",  x"6c",  x"0d",  x"66",  x"6c",  x"f8",  x"bc", -- 31A8
         x"00",  x"62",  x"68",  x"78",  x"68",  x"25",  x"62",  x"fe", -- 31B0
         x"07",  x"24",  x"60",  x"f0",  x"1f",  x"57",  x"ce",  x"1f", -- 31B8
         x"32",  x"7a",  x"36",  x"37",  x"78",  x"41",  x"c0",  x"ce", -- 31C0
         x"47",  x"1e",  x"0c",  x"00",  x"c1",  x"8f",  x"e6",  x"b1", -- 31C8
         x"34",  x"70",  x"3a",  x"e6",  x"00",  x"f0",  x"42",  x"9e", -- 31D0
         x"62",  x"60",  x"66",  x"37",  x"c6",  x"ee",  x"fe",  x"d6", -- 31D8
         x"c6",  x"f0",  x"00",  x"07",  x"e6",  x"f6",  x"de",  x"ce", -- 31E0
         x"58",  x"c6",  x"c7",  x"d6",  x"0d",  x"cb",  x"32",  x"7f", -- 31E8
         x"6f",  x"21",  x"4f",  x"7e",  x"89",  x"00",  x"dc",  x"78", -- 31F0
         x"1c",  x"2f",  x"0f",  x"37",  x"97",  x"00",  x"f0",  x"3c", -- 31F8
         x"0e",  x"c6",  x"69",  x"7c",  x"0f",  x"b4",  x"7b",  x"57", -- 3200
         x"1d",  x"00",  x"be",  x"07",  x"04",  x"bc",  x"6b",  x"47", -- 3208
         x"00",  x"d6",  x"fe",  x"77",  x"ee",  x"47",  x"44",  x"52", -- 3210
         x"4a",  x"58",  x"17",  x"27",  x"fe",  x"c6",  x"8c",  x"29", -- 3218
         x"18",  x"32",  x"6f",  x"ff",  x"32",  x"00",  x"18",  x"5a", -- 3220
         x"00",  x"fd",  x"12",  x"06",  x"06",  x"c5",  x"fa",  x"10", -- 3228
         x"f1",  x"2d",  x"2c",  x"23",  x"00",  x"ff",  x"c3",  x"bf", -- 3230
         x"aa",  x"36",  x"47",  x"02",  x"63",  x"db",  x"02",  x"77", -- 3238
         x"02",  x"33",  x"02",  x"6d",  x"b0",  x"02",  x"f6",  x"02", -- 3240
         x"27",  x"b5",  x"02",  x"7a",  x"02",  x"99",  x"66",  x"94", -- 3248
         x"06",  x"cd",  x"c9",  x"1b",  x"18",  x"07",  x"37",  x"08", -- 3250
         x"21",  x"cd",  x"12",  x"c8",  x"c0",  x"f5",  x"db",  x"88", -- 3258
         x"05",  x"cb",  x"d7",  x"d3",  x"88",  x"f1",  x"5a",  x"0f", -- 3260
         x"0a",  x"97",  x"8f",  x"0a",  x"c9",  x"f3",  x"ed",  x"94", -- 3268
         x"e1",  x"df",  x"c0",  x"3b",  x"3b",  x"fb",  x"f5",  x"d5", -- 3270
         x"00",  x"5e",  x"16",  x"00",  x"2a",  x"b0",  x"b7",  x"19", -- 3278
         x"19",  x"a7",  x"a7",  x"f4",  x"e1",  x"f1",  x"e3",  x"29", -- 3280
         x"c9",  x"a7",  x"a2",  x"f4",  x"ea",  x"0f",  x"bb",  x"f0", -- 3288
         x"e3",  x"e5",  x"1b",  x"f3",  x"a0",  x"3a",  x"80",  x"b7", -- 3290
         x"5f",  x"00",  x"18",  x"dd",  x"37",  x"18",  x"ea",  x"c1", -- 3298
         x"fd",  x"e5",  x"55",  x"fd",  x"c7",  x"01",  x"fd",  x"39", -- 32A0
         x"f3",  x"dd",  x"77",  x"0b",  x"66",  x"52",  x"cb",  x"ef", -- 32A8
         x"49",  x"ed",  x"03",  x"7b",  x"ae",  x"b7",  x"fb",  x"dd", -- 32B0
         x"7e",  x"ed",  x"8d",  x"83",  x"65",  x"15",  x"0c",  x"97", -- 32B8
         x"cb",  x"af",  x"f3",  x"16",  x"fd",  x"f9",  x"b3",  x"14", -- 32C0
         x"fd",  x"e1",  x"16",  x"50",  x"e3",  x"55",  x"23",  x"eb", -- 32C8
         x"19",  x"1b",  x"eb",  x"e3",  x"d5",  x"21",  x"d1",  x"d0", -- 32D0
         x"50",  x"31",  x"c4",  x"01",  x"af",  x"1b",  x"47",  x"4f", -- 32D8
         x"02",  x"eb",  x"80",  x"fc",  x"10",  x"fa",  x"0e",  x"80", -- 32E0
         x"ed",  x"79",  x"00",  x"10",  x"fc",  x"cd",  x"d0",  x"f3", -- 32E8
         x"af",  x"32",  x"9b",  x"d4",  x"86",  x"bb",  x"f6",  x"7a", -- 32F0
         x"3c",  x"c8",  x"38",  x"df",  x"af",  x"ff",  x"46",  x"3e", -- 32F8
         x"cb",  x"ee",  x"29",  x"f8",  x"35",  x"8b",  x"06",  x"cd", -- 3300
         x"61",  x"fb",  x"cd",  x"d9",  x"ad",  x"c1",  x"6d",  x"fb", -- 3308
         x"18",  x"06",  x"54",  x"36",  x"27",  x"3a",  x"36",  x"00", -- 3310
         x"a8",  x"e1",  x"5b",  x"0c",  x"16",  x"d5",  x"d2",  x"a5", -- 3318
         x"c3",  x"83",  x"19",  x"01",  x"80",  x"08",  x"ed",  x"78", -- 3320
         x"13",  x"18",  x"1c",  x"3e",  x"43",  x"4a",  x"32",  x"08", -- 3328
         x"b8",  x"c6",  x"73",  x"04",  x"e6",  x"fc",  x"87",  x"00", -- 3330
         x"04",  x"d3",  x"86",  x"c3",  x"00",  x"01",  x"40",  x"7f", -- 3338
         x"7f",  x"4d",  x"45",  x"4e",  x"55",  x"c0",  x"a9",  x"cd", -- 3340
         x"ee",  x"f1",  x"7e",  x"0c",  x"e6",  x"20",  x"00",  x"4b", -- 3348
         x"43",  x"2d",  x"43",  x"41",  x"4f",  x"53",  x"20",  x"03", -- 3350
         x"34",  x"2e",  x"32",  x"20",  x"2a",  x"00",  x"c8",  x"06", -- 3358
         x"c0",  x"1d",  x"cd",  x"28",  x"6b",  x"f3",  x"1c",  x"02", -- 3360
         x"25",  x"f8",  x"a7",  x"de",  x"e3",  x"30",  x"38",  x"29", -- 3368
         x"3c",  x"09",  x"ed",  x"b1",  x"e2",  x"03",  x"83",  x"f1", -- 3370
         x"ed",  x"a1",  x"20",  x"f7",  x"df",  x"70",  x"02",  x"38", -- 3378
         x"e1",  x"fe",  x"0c",  x"30",  x"38",  x"e0",  x"fe",  x"ff", -- 3380
         x"c0",  x"dc",  x"cd",  x"1d",  x"f2",  x"23",  x"0b",  x"ff", -- 3388
         x"fd",  x"48",  x"5d",  x"61",  x"2e",  x"07",  x"2d",  x"34", -- 3390
         x"f3",  x"13",  x"1a",  x"8a",  x"87",  x"28",  x"f2",  x"ef", -- 3398
         x"00",  x"ef",  x"cd",  x"a9",  x"f1",  x"30",  x"72",  x"e7", -- 33A0
         x"e9",  x"c7",  x"66",  x"f3",  x"2a",  x"21",  x"7e",  x"bb", -- 33A8
         x"3b",  x"e4",  x"ec",  x"f3",  x"cd",  x"02",  x"eb",  x"f4", -- 33B0
         x"c0",  x"c3",  x"3e",  x"f0",  x"89",  x"61",  x"45",  x"4d", -- 33B8
         x"05",  x"53",  x"37",  x"3f",  x"e0",  x"e2",  x"53",  x"cc", -- 33C0
         x"1a",  x"06",  x"13",  x"fe",  x"21",  x"38",  x"08",  x"0b", -- 33C8
         x"28",  x"63",  x"f6",  x"e6",  x"bd",  x"b0",  x"b0",  x"63", -- 33D0
         x"07",  x"46",  x"38",  x"f3",  x"23",  x"18",  x"00",  x"f4", -- 33D8
         x"f1",  x"f1",  x"37",  x"c9",  x"3d",  x"c8",  x"f5",  x"ce", -- 33E0
         x"15",  x"fa",  x"47",  x"8e",  x"01",  x"da",  x"f1",  x"10", -- 33E8
         x"fb",  x"c9",  x"85",  x"39",  x"02",  x"cd",  x"76",  x"f3", -- 33F0
         x"05",  x"50",  x"a7",  x"ca",  x"61",  x"f0",  x"03",  x"81", -- 33F8
         x"18",  x"99",  x"13",  x"0a",  x"f2",  x"8c",  x"c0",  x"fb", -- 3400
         x"e5",  x"2a",  x"b9",  x"1e",  x"b7",  x"e3",  x"22",  x"03", -- 3408
         x"ca",  x"25",  x"21",  x"a4",  x"2b",  x"0c",  x"bb",  x"0c", -- 3410
         x"03",  x"ec",  x"0c",  x"09",  x"18",  x"04",  x"bc",  x"1c", -- 3418
         x"bb",  x"a5",  x"cf",  x"26",  x"f5",  x"d0",  x"4b",  x"f1", -- 3420
         x"d1",  x"2c",  x"82",  x"d6",  x"e1",  x"f8",  x"34",  x"d3", -- 3428
         x"40",  x"dd",  x"cb",  x"08",  x"76",  x"20",  x"4c",  x"76", -- 3430
         x"f3",  x"ee",  x"af",  x"d1",  x"80",  x"13",  x"5f",  x"cd", -- 3438
         x"4a",  x"f7",  x"1c",  x"31",  x"06",  x"0f",  x"cd",  x"c0", -- 3440
         x"fd",  x"1b",  x"0b",  x"00",  x"78",  x"b1",  x"20",  x"f6", -- 3448
         x"18",  x"ee",  x"cd",  x"40",  x"00",  x"e0",  x"cb",  x"cd", -- 3450
         x"cb",  x"d5",  x"7e",  x"47",  x"ee",  x"28",  x"7f",  x"77", -- 3458
         x"17",  x"30",  x"fb",  x"03",  x"70",  x"18",  x"05",  x"cb", -- 3460
         x"43",  x"c4",  x"27",  x"51",  x"57",  x"3d",  x"6e",  x"01", -- 3468
         x"c8",  x"dc",  x"c4",  x"05",  x"e3",  x"00",  x"7a",  x"21", -- 3470
         x"a2",  x"b7",  x"cb",  x"66",  x"28",  x"0d",  x"90",  x"49", -- 3478
         x"63",  x"e1",  x"30",  x"ed",  x"53",  x"06",  x"18",  x"a9", -- 3480
         x"fe",  x"1b",  x"00",  x"20",  x"04",  x"cb",  x"e6",  x"18", -- 3488
         x"a1",  x"fe",  x"f1",  x"2b",  x"38",  x"90",  x"2a",  x"a2", -- 3490
         x"77",  x"0f",  x"f1",  x"01",  x"00",  x"b9",  x"7e",  x"a7", -- 3498
         x"d0",  x"a7",  x"fb",  x"10",  x"f9",  x"2c",  x"18",  x"08", -- 34A0
         x"e1",  x"41",  x"1b",  x"2a",  x"d1",  x"b7",  x"7e",  x"5d", -- 34A8
         x"27",  x"df",  x"3b",  x"22",  x"08",  x"43",  x"0b",  x"e6", -- 34B0
         x"c3",  x"3b",  x"f2",  x"0b",  x"14",  x"a7",  x"20",  x"07", -- 34B8
         x"32",  x"b6",  x"12",  x"c3",  x"41",  x"f2",  x"08",  x"59", -- 34C0
         x"ca",  x"34",  x"f2",  x"aa",  x"5a",  x"23",  x"29",  x"22", -- 34C8
         x"e3",  x"f9",  x"3f",  x"bb",  x"a0",  x"04",  x"39",  x"60", -- 34D0
         x"e2",  x"00",  x"6b",  x"ee",  x"9a",  x"79",  x"03",  x"91", -- 34D8
         x"86",  x"a8",  x"fb",  x"c8",  x"fc",  x"ea",  x"63",  x"c3", -- 34E0
         x"12",  x"f0",  x"95",  x"1c",  x"8a",  x"44",  x"c3",  x"53", -- 34E8
         x"f3",  x"40",  x"02",  x"82",  x"dc",  x"00",  x"03",  x"b2", -- 34F0
         x"db",  x"ed",  x"0b",  x"05",  x"00",  x"22",  x"00",  x"08", -- 34F8
         x"09",  x"a8",  x"09",  x"06",  x"cd",  x"17",  x"f2",  x"a1", -- 3500
         x"c1",  x"f3",  x"9a",  x"e0",  x"0a",  x"f1",  x"2b",  x"5a", -- 3508
         x"60",  x"ba",  x"ab",  x"3a",  x"f8",  x"f9",  x"57",  x"15", -- 3510
         x"50",  x"e5",  x"88",  x"b1",  x"eb",  x"9b",  x"50",  x"7c", -- 3518
         x"e9",  x"a8",  x"7d",  x"03",  x"3e",  x"20",  x"74",  x"c3", -- 3520
         x"26",  x"e2",  x"40",  x"45",  x"52",  x"52",  x"4f",  x"52", -- 3528
         x"28",  x"07",  x"00",  x"09",  x"0d",  x"0a",  x"00",  x"00", -- 3530
         x"c9",  x"3e",  x"10",  x"18",  x"e8",  x"f5",  x"1f",  x"a0", -- 3538
         x"00",  x"cd",  x"7f",  x"f3",  x"f1",  x"c0",  x"d6",  x"c6", -- 3540
         x"90",  x"07",  x"27",  x"ce",  x"40",  x"27",  x"18",  x"df", -- 3548
         x"4c",  x"8c",  x"8d",  x"c2",  x"54",  x"f3",  x"eb",  x"c9", -- 3550
         x"43",  x"8a",  x"01",  x"fa",  x"af",  x"21",  x"98",  x"b7", -- 3558
         x"77",  x"2b",  x"43",  x"01",  x"1a",  x"b7",  x"c8",  x"0f", -- 3560
         x"0a",  x"c8",  x"d6",  x"30",  x"d8",  x"cc",  x"40",  x"0b", -- 3568
         x"d6",  x"07",  x"e6",  x"78",  x"df",  x"07",  x"0a",  x"10", -- 3570
         x"3f",  x"d8",  x"05",  x"13",  x"34",  x"23",  x"ed",  x"6f", -- 3578
         x"03",  x"02",  x"2b",  x"2b",  x"28",  x"dc",  x"1b",  x"ec", -- 3580
         x"2b",  x"c4",  x"41",  x"0e",  x"c7",  x"c3",  x"a1",  x"c1", -- 3588
         x"11",  x"99",  x"88",  x"8a",  x"f4",  x"f2",  x"01",  x"07", -- 3590
         x"34",  x"00",  x"ed",  x"b0",  x"0e",  x"b6",  x"2d",  x"dd", -- 3598
         x"05",  x"21",  x"d8",  x"ef",  x"22",  x"00",  x"b8",  x"c4", -- 35A0
         x"bb",  x"03",  x"22",  x"01",  x"02",  x"b8",  x"3e",  x"03", -- 35A8
         x"32",  x"04",  x"b8",  x"86",  x"b1",  x"d0",  x"40",  x"07", -- 35B0
         x"21",  x"63",  x"f4",  x"cd",  x"00",  x"5a",  x"f4",  x"dd", -- 35B8
         x"21",  x"f0",  x"01",  x"dd",  x"36",  x"33",  x"01",  x"28", -- 35C0
         x"03",  x"04",  x"63",  x"c3",  x"b0",  x"21",  x"ba",  x"fc", -- 35C8
         x"32",  x"01",  x"d7",  x"b7",  x"1e",  x"e2",  x"57",  x"01", -- 35D0
         x"0e",  x"46",  x"3d",  x"dd",  x"66",  x"1a",  x"6e",  x"56", -- 35D8
         x"04",  x"ca",  x"61",  x"1c",  x"08",  x"88",  x"dd",  x"74", -- 35E0
         x"99",  x"0c",  x"75",  x"04",  x"09",  x"0e",  x"3a",  x"99", -- 35E8
         x"03",  x"0f",  x"fc",  x"03",  x"09",  x"7f",  x"4c",  x"45", -- 35F0
         x"3a",  x"2c",  x"ed",  x"47",  x"0b",  x"16",  x"04",  x"21", -- 35F8
         x"7b",  x"4a",  x"f1",  x"13",  x"9e",  x"c3",  x"03",  x"06", -- 3600
         x"b7",  x"c9",  x"c5",  x"86",  x"f6",  x"46",  x"97",  x"0d", -- 3608
         x"b3",  x"a6",  x"f0",  x"ce",  x"06",  x"51",  x"f4",  x"15", -- 3610
         x"20",  x"fa",  x"fa",  x"60",  x"8a",  x"01",  x"e4",  x"88", -- 3618
         x"01",  x"03",  x"0f",  x"8a",  x"02",  x"0f",  x"03",  x"8b", -- 3620
         x"90",  x"d0",  x"0f",  x"83",  x"89",  x"01",  x"31",  x"ff", -- 3628
         x"84",  x"72",  x"86",  x"01",  x"63",  x"40",  x"17",  x"8b", -- 3630
         x"01",  x"e6",  x"8c",  x"01",  x"06",  x"e8",  x"8e",  x"02", -- 3638
         x"47",  x"0c",  x"dd",  x"a0",  x"53",  x"41",  x"56",  x"45", -- 3640
         x"01",  x"d1",  x"c3",  x"da",  x"22",  x"95",  x"9a",  x"4e", -- 3648
         x"41",  x"ce",  x"96",  x"20",  x"3a",  x"9a",  x"ae",  x"21", -- 3650
         x"b6",  x"00",  x"19",  x"11",  x"00",  x"b7",  x"01",  x"0b", -- 3658
         x"a0",  x"93",  x"0c",  x"af",  x"12",  x"21",  x"81",  x"a0", -- 3660
         x"06",  x"10",  x"0e",  x"15",  x"0a",  x"cd",  x"6d",  x"48", -- 3668
         x"75",  x"1c",  x"9f",  x"3d",  x"c0",  x"c1",  x"97",  x"05", -- 3670
         x"82",  x"9d",  x"06",  x"d7",  x"f7",  x"2d",  x"32",  x"e8", -- 3678
         x"f1",  x"a2",  x"5a",  x"a0",  x"fd",  x"83",  x"da",  x"e0", -- 3680
         x"e4",  x"11",  x"80",  x"37",  x"c9",  x"9b",  x"84",  x"80", -- 3688
         x"a2",  x"52",  x"d2",  x"d9",  x"00",  x"e4",  x"cd",  x"2b", -- 3690
         x"e5",  x"18",  x"d6",  x"ed",  x"4b",  x"2e",  x"86",  x"b7", -- 3698
         x"11",  x"9e",  x"34",  x"3a",  x"46",  x"91",  x"af",  x"34", -- 36A0
         x"93",  x"82",  x"91",  x"e5",  x"30",  x"20",  x"9a",  x"3a", -- 36A8
         x"09",  x"00",  x"20",  x"ce",  x"3d",  x"20",  x"3f",  x"e8", -- 36B0
         x"f5",  x"a8",  x"03",  x"03",  x"3d",  x"28",  x"e6",  x"cd", -- 36B8
         x"38",  x"df",  x"23",  x"03",  x"37",  x"fa",  x"11",  x"0a", -- 36C0
         x"20",  x"db",  x"4a",  x"b9",  x"dd",  x"3e",  x"46",  x"03", -- 36C8
         x"9d",  x"62",  x"17",  x"ba",  x"28",  x"0a",  x"0b",  x"3c", -- 36D0
         x"28",  x"08",  x"27",  x"3c",  x"2a",  x"19",  x"f7",  x"56", -- 36D8
         x"c3",  x"07",  x"e0",  x"5e",  x"08",  x"e7",  x"a5",  x"20", -- 36E0
         x"ed",  x"1e",  x"86",  x"e0",  x"23",  x"b7",  x"06",  x"0b", -- 36E8
         x"dd",  x"5a",  x"e9",  x"7d",  x"9e",  x"0b",  x"c3",  x"5c", -- 36F0
         x"c2",  x"06",  x"3f",  x"00",  x"00",  x"61",  x"c3",  x"87", -- 36F8
         x"86",  x"d8",  x"d6",  x"01",  x"52",  x"49",  x"46",  x"59", -- 3700
         x"88",  x"c0",  x"cb",  x"07",  x"86",  x"30",  x"18",  x"0b", -- 3708
         x"0e",  x"4c",  x"4f",  x"41",  x"44",  x"bd",  x"0c",  x"ef", -- 3710
         x"ca",  x"b4",  x"e4",  x"c5",  x"0c",  x"b4",  x"58",  x"03", -- 3718
         x"7a",  x"fa",  x"f4",  x"38",  x"50",  x"d4",  x"12",  x"46", -- 3720
         x"28",  x"49",  x"3c",  x"2e",  x"10",  x"6f",  x"e5",  x"9b", -- 3728
         x"e3",  x"f4",  x"86",  x"07",  x"7e",  x"cb",  x"27",  x"01", -- 3730
         x"e6",  x"0b",  x"1c",  x"dd",  x"b6",  x"07",  x"0c",  x"03", -- 3738
         x"d6",  x"02",  x"fe",  x"09",  x"30",  x"a9",  x"c2",  x"05", -- 3740
         x"15",  x"03",  x"c2",  x"13",  x"c2",  x"05",  x"11",  x"86", -- 3748
         x"c2",  x"af",  x"e7",  x"13",  x"c5",  x"11",  x"81",  x"cd", -- 3750
         x"09",  x"eb",  x"d0",  x"01",  x"3d",  x"66",  x"20",  x"03", -- 3758
         x"03",  x"e3",  x"09",  x"e3",  x"c1",  x"ed",  x"43",  x"e2", -- 3760
         x"01",  x"cd",  x"89",  x"f3",  x"40",  x"93",  x"eb",  x"b4", -- 3768
         x"57",  x"a6",  x"86",  x"57",  x"12",  x"e5",  x"87",  x"3c", -- 3770
         x"dc",  x"62",  x"c2",  x"42",  x"ca",  x"44",  x"01",  x"4d", -- 3778
         x"ab",  x"0c",  x"c0",  x"72",  x"d7",  x"06",  x"34",  x"02", -- 3780
         x"20",  x"de",  x"cd",  x"a0",  x"17",  x"6f",  x"82",  x"f2", -- 3788
         x"c0",  x"de",  x"06",  x"1c",  x"e9",  x"e1",  x"8e",  x"a1", -- 3790
         x"a8",  x"d8",  x"2a",  x"b0",  x"41",  x"e9",  x"a8",  x"30", -- 3798
         x"43",  x"4f",  x"aa",  x"ec",  x"34",  x"d9",  x"ca",  x"63", -- 37A0
         x"c1",  x"d9",  x"35",  x"e5",  x"af",  x"cc",  x"30",  x"a1", -- 37A8
         x"d1",  x"cb",  x"9e",  x"a6",  x"e2",  x"1d",  x"44",  x"02", -- 37B0
         x"49",  x"53",  x"50",  x"4c",  x"41",  x"59",  x"42",  x"1f", -- 37B8
         x"42",  x"c2",  x"aa",  x"1f",  x"be",  x"4e",  x"7e",  x"c3", -- 37C0
         x"0c",  x"a5",  x"a6",  x"4f",  x"a5",  x"1b",  x"46",  x"18", -- 37C8
         x"0a",  x"6a",  x"c2",  x"18",  x"e5",  x"17",  x"18",  x"77", -- 37D0
         x"18",  x"e6",  x"16",  x"57",  x"49",  x"4e",  x"33",  x"44", -- 37D8
         x"4f",  x"db",  x"c1",  x"b4",  x"2a",  x"88",  x"df",  x"26", -- 37E0
         x"65",  x"69",  x"1d",  x"53",  x"3a",  x"88",  x"88",  x"d0", -- 37E8
         x"c4",  x"00",  x"fe",  x"04",  x"20",  x"05",  x"38",  x"09", -- 37F0
         x"af",  x"0c",  x"18",  x"03",  x"3a",  x"8a",  x"b6",  x"0a", -- 37F8
         x"94",  x"f6",  x"fe",  x"29",  x"11",  x"cc",  x"2d",  x"6a", -- 3800
         x"72",  x"7d",  x"c5",  x"ab",  x"cb",  x"a0",  x"ae",  x"f6", -- 3808
         x"d8",  x"eb",  x"37",  x"11",  x"9c",  x"95",  x"30",  x"1b", -- 3810
         x"c6",  x"08",  x"87",  x"5f",  x"87",  x"87",  x"07",  x"83", -- 3818
         x"5f",  x"16",  x"b9",  x"a7",  x"87",  x"8b",  x"3a",  x"1a", -- 3820
         x"c3",  x"31",  x"5b",  x"e0",  x"f1",  x"21",  x"1c",  x"28", -- 3828
         x"01",  x"0a",  x"a0",  x"cd",  x"c9",  x"23",  x"a1",  x"c6", -- 3830
         x"c8",  x"cd",  x"2a",  x"f8",  x"ec",  x"f7",  x"6f",  x"4b", -- 3838
         x"45",  x"c0",  x"83",  x"fe",  x"01",  x"3d",  x"c0",  x"7d", -- 3840
         x"10",  x"a9",  x"92",  x"d0",  x"3f",  x"bc",  x"fb",  x"16", -- 3848
         x"bc",  x"fd",  x"f8",  x"05",  x"f6",  x"f5",  x"2b",  x"f1", -- 3850
         x"30",  x"c3",  x"fe",  x"13",  x"ca",  x"c5",  x"a3",  x"f5", -- 3858
         x"9e",  x"de",  x"c0",  x"4c",  x"15",  x"35",  x"28",  x"ed", -- 3860
         x"00",  x"54",  x"5d",  x"e5",  x"23",  x"3e",  x"9c",  x"95", -- 3868
         x"4f",  x"a1",  x"9a",  x"5c",  x"f1",  x"a0",  x"8c",  x"da", -- 3870
         x"3a",  x"9a",  x"64",  x"20",  x"d6",  x"1b",  x"e5",  x"3e", -- 3878
         x"9b",  x"13",  x"21",  x"0a",  x"06",  x"11",  x"9b",  x"b9", -- 3880
         x"ed",  x"b8",  x"19",  x"23",  x"5a",  x"77",  x"5e",  x"c1", -- 3888
         x"46",  x"5e",  x"4c",  x"82",  x"29",  x"54",  x"00",  x"e6", -- 3890
         x"f7",  x"c0",  x"a0",  x"ac",  x"15",  x"d5",  x"f5",  x"e5", -- 3898
         x"ed",  x"00",  x"38",  x"0a",  x"c5",  x"06",  x"08",  x"0f", -- 38A0
         x"7e",  x"2f",  x"77",  x"2c",  x"8f",  x"1a",  x"c1",  x"2d", -- 38A8
         x"d1",  x"e4",  x"a7",  x"a7",  x"f5",  x"28",  x"2a",  x"d3", -- 38B0
         x"b5",  x"8e",  x"d5",  x"b7",  x"c7",  x"45",  x"c3",  x"ec", -- 38B8
         x"f7",  x"ac",  x"2f",  x"e4",  x"dc",  x"1a",  x"3a",  x"8d", -- 38C0
         x"0c",  x"4f",  x"69",  x"af",  x"2c",  x"cb",  x"1d",  x"c8", -- 38C8
         x"92",  x"81",  x"1f",  x"c6",  x"05",  x"10",  x"f8",  x"67", -- 38D0
         x"82",  x"00",  x"79",  x"cb",  x"21",  x"cb",  x"10",  x"f0", -- 38D8
         x"fd",  x"01",  x"01",  x"18",  x"00",  x"d9",  x"4f",  x"99", -- 38E0
         x"1e",  x"cd",  x"c2",  x"2e",  x"02",  x"d9",  x"64",  x"a7", -- 38E8
         x"b6",  x"03",  x"64",  x"03",  x"bf",  x"19",  x"03",  x"d9", -- 38F0
         x"30",  x"0c",  x"d9",  x"e3",  x"eb",  x"0d",  x"1e",  x"52", -- 38F8
         x"1b",  x"1b",  x"ff",  x"00",  x"d9",  x"0d",  x"04",  x"79", -- 3900
         x"b8",  x"30",  x"dd",  x"f5",  x"fa",  x"78",  x"e1",  x"85", -- 3908
         x"af",  x"57",  x"44",  x"b1",  x"e5",  x"06",  x"59",  x"19", -- 3910
         x"cd",  x"d6",  x"f7",  x"0a",  x"e1",  x"76",  x"59",  x"20", -- 3918
         x"98",  x"aa",  x"58",  x"28",  x"68",  x"d1",  x"a4",  x"f7", -- 3920
         x"1d",  x"d5",  x"57",  x"58",  x"ba",  x"28",  x"d1",  x"87", -- 3928
         x"06",  x"f5",  x"7d",  x"e6",  x"f4",  x"6c",  x"f8",  x"56", -- 3930
         x"fd",  x"7d",  x"12",  x"cb",  x"3c",  x"1f",  x"80",  x"02", -- 3938
         x"fe",  x"28",  x"30",  x"31",  x"f6",  x"80",  x"67",  x"1e", -- 3940
         x"3e",  x"ff",  x"82",  x"af",  x"07",  x"ab",  x"6f",  x"3a", -- 3948
         x"d6",  x"c3",  x"0c",  x"0a",  x"ae",  x"c0",  x"01",  x"5e", -- 3950
         x"28",  x"2d",  x"cb",  x"4a",  x"0d",  x"20",  x"23",  x"cb", -- 3958
         x"42",  x"de",  x"0c",  x"b6",  x"77",  x"97",  x"c3",  x"01", -- 3960
         x"5f",  x"ee",  x"02",  x"83",  x"e3",  x"84",  x"7e",  x"3d", -- 3968
         x"19",  x"b2",  x"77",  x"7b",  x"07",  x"fb",  x"f1",  x"74", -- 3970
         x"ff",  x"ae",  x"00",  x"cb",  x"82",  x"c3",  x"20",  x"f8", -- 3978
         x"2f",  x"a6",  x"77",  x"fc",  x"b4",  x"f8",  x"47",  x"0e", -- 3980
         x"b6",  x"cb",  x"5a",  x"20",  x"9b",  x"6d",  x"2a",  x"4f", -- 3988
         x"23",  x"2a",  x"78",  x"10",  x"5a",  x"62",  x"10",  x"79", -- 3990
         x"8b",  x"2d",  x"18",  x"d0",  x"f1",  x"00",  x"7c",  x"c1", -- 3998
         x"18",  x"28",  x"b0",  x"07",  x"2b",  x"c7",  x"18",  x"20", -- 39A0
         x"b6",  x"07",  x"a7",  x"07",  x"18",  x"a3",  x"98",  x"15", -- 39A8
         x"2a",  x"c9",  x"b7",  x"d2",  x"e9",  x"e9",  x"0c",  x"b3", -- 39B0
         x"55",  x"4c",  x"90",  x"cb",  x"56",  x"00",  x"cb",  x"34", -- 39B8
         x"8d",  x"ec",  x"59",  x"db",  x"7c",  x"ef",  x"90",  x"11", -- 39C0
         x"28",  x"c0",  x"f4",  x"ac",  x"e5",  x"c5",  x"00",  x"cd", -- 39C8
         x"7a",  x"f0",  x"cb",  x"6b",  x"d5",  x"20",  x"53",  x"60", -- 39D0
         x"23",  x"97",  x"7b",  x"0c",  x"20",  x"42",  x"e5",  x"7b", -- 39D8
         x"8d",  x"00",  x"21",  x"f1",  x"f8",  x"85",  x"6f",  x"7a", -- 39E0
         x"3d",  x"53",  x"5e",  x"c8",  x"0f",  x"77",  x"f0",  x"d1", -- 39E8
         x"57",  x"10",  x"7b",  x"3d",  x"43",  x"20",  x"54",  x"f8", -- 39F0
         x"65",  x"ef",  x"5d",  x"cb",  x"86",  x"28",  x"59",  x"29", -- 39F8
         x"c1",  x"f6",  x"c8",  x"c0",  x"59",  x"cc",  x"6a",  x"f5", -- 3A00
         x"7a",  x"2b",  x"cb",  x"9b",  x"69",  x"92",  x"20",  x"c9", -- 3A08
         x"16",  x"24",  x"37",  x"1d",  x"38",  x"06",  x"02",  x"f8", -- 3A10
         x"8c",  x"cd",  x"ca",  x"e3",  x"34",  x"30",  x"e8",  x"01", -- 3A18
         x"cb",  x"bb",  x"18",  x"e4",  x"3a",  x"5e",  x"03",  x"92", -- 3A20
         x"ff",  x"09",  x"85",  x"1e",  x"cd",  x"41",  x"c6",  x"7e", -- 3A28
         x"66",  x"f5",  x"e6",  x"55",  x"5f",  x"87",  x"fb",  x"fe", -- 3A30
         x"46",  x"b0",  x"c8",  x"b3",  x"89",  x"57",  x"f7",  x"82", -- 3A38
         x"55",  x"d0",  x"b8",  x"4e",  x"cc",  x"1c",  x"c5",  x"0e", -- 3A40
         x"8c",  x"eb",  x"0a",  x"f9",  x"0c",  x"eb",  x"04",  x"00", -- 3A48
         x"c1",  x"79",  x"ee",  x"1f",  x"f6",  x"81",  x"4f",  x"78", -- 3A50
         x"c5",  x"39",  x"0d",  x"cb",  x"b9",  x"01",  x"1d",  x"ce", -- 3A58
         x"3e",  x"c7",  x"d3",  x"8e",  x"78",  x"80",  x"02",  x"06", -- 3A60
         x"60",  x"db",  x"89",  x"a0",  x"b1",  x"d3",  x"33",  x"89", -- 3A68
         x"c9",  x"f8",  x"37",  x"2e",  x"03",  x"b0",  x"00",  x"6f", -- 3A70
         x"3e",  x"07",  x"cb",  x"44",  x"28",  x"02",  x"f6",  x"dc", -- 3A78
         x"a4",  x"79",  x"ed",  x"7b",  x"69",  x"e3",  x"d8",  x"c8", -- 3A80
         x"22",  x"cb",  x"b7",  x"a1",  x"a7",  x"31",  x"e6",  x"f8", -- 3A88
         x"9a",  x"d9",  x"d6",  x"01",  x"49",  x"10",  x"ad",  x"42", -- 3A90
         x"10",  x"f6",  x"05",  x"18",  x"ed",  x"7c",  x"0c",  x"1d", -- 3A98
         x"fe",  x"f6",  x"13",  x"04",  x"18",  x"de",  x"ff",  x"2c", -- 3AA0
         x"1b",  x"10",  x"f2",  x"8a",  x"cf",  x"fe",  x"50",  x"7e", -- 3AA8
         x"ee",  x"04",  x"77",  x"56",  x"c9",  x"10",  x"e4",  x"26", -- 3AB0
         x"18",  x"c0",  x"65",  x"ee",  x"76",  x"80",  x"65",  x"0c", -- 3AB8
         x"08",  x"29",  x"18",  x"b3",  x"e4",  x"c2",  x"32",  x"34", -- 3AC0
         x"4f",  x"55",  x"54",  x"8d",  x"00",  x"d5",  x"c2",  x"3e", -- 3AC8
         x"0d",  x"cd",  x"06",  x"fa",  x"3e",  x"55",  x"0a",  x"04", -- 3AD0
         x"b5",  x"97",  x"1f",  x"12",  x"cf",  x"c3",  x"ef",  x"49", -- 3AD8
         x"23",  x"8a",  x"e5",  x"50",  x"43",  x"23",  x"4f",  x"c6", -- 3AE0
         x"f6",  x"0b",  x"07",  x"6a",  x"c3",  x"07",  x"dc",  x"b3", -- 3AE8
         x"8d",  x"ca",  x"5b",  x"e1",  x"db",  x"00",  x"7f",  x"28", -- 3AF0
         x"29",  x"e6",  x"f0",  x"fe",  x"90",  x"e0",  x"e8",  x"fe", -- 3AF8
         x"a0",  x"18",  x"20",  x"1f",  x"f1",  x"f1",  x"8f",  x"21", -- 3B00
         x"92",  x"fb",  x"a0",  x"b5",  x"d4",  x"f8",  x"c7",  x"0f", -- 3B08
         x"0e",  x"00",  x"06",  x"09",  x"7e",  x"18",  x"09",  x"f1", -- 3B10
         x"fe",  x"7e",  x"0f",  x"20",  x"08",  x"3e",  x"83",  x"96", -- 3B18
         x"f1",  x"c5",  x"6c",  x"f5",  x"0b",  x"09",  x"f7",  x"3a", -- 3B20
         x"35",  x"91",  x"71",  x"5f",  x"28",  x"0e",  x"8e",  x"0c", -- 3B28
         x"7f",  x"20",  x"02",  x"8b",  x"7c",  x"a7",  x"66",  x"30", -- 3B30
         x"05",  x"5f",  x"f5",  x"a9",  x"4a",  x"d4",  x"7b",  x"c4", -- 3B38
         x"99",  x"ed",  x"78",  x"2b",  x"cb",  x"57",  x"2f",  x"6e", -- 3B40
         x"db",  x"9e",  x"fc",  x"21",  x"ea",  x"c1",  x"f1",  x"9d", -- 3B48
         x"ff",  x"b6",  x"18",  x"08",  x"18",  x"f1",  x"8a",  x"3d", -- 3B50
         x"9d",  x"d2",  x"26",  x"e1",  x"17",  x"26",  x"c6",  x"18", -- 3B58
         x"18",  x"d7",  x"c5",  x"b0",  x"94",  x"07",  x"c5",  x"99", -- 3B60
         x"21",  x"47",  x"b1",  x"a2",  x"3e",  x"05",  x"9c",  x"36", -- 3B68
         x"3e",  x"ea",  x"03",  x"8b",  x"0d",  x"07",  x"ff",  x"e1", -- 3B70
         x"15",  x"18",  x"f3",  x"22",  x"14",  x"6a",  x"af",  x"4f", -- 3B78
         x"57",  x"19",  x"d3",  x"97",  x"58",  x"d6",  x"44",  x"f9", -- 3B80
         x"cd",  x"19",  x"54",  x"0e",  x"01",  x"a3",  x"82",  x"0d", -- 3B88
         x"9e",  x"5d",  x"0c",  x"e8",  x"ba",  x"b8",  x"f1",  x"d0", -- 3B90
         x"fe",  x"db",  x"09",  x"07",  x"f5",  x"3e",  x"18",  x"d3", -- 3B98
         x"0b",  x"33",  x"fe",  x"03",  x"33",  x"03",  x"e4",  x"c6", -- 3BA0
         x"57",  x"fb",  x"99",  x"e7",  x"28",  x"0a",  x"c1",  x"fc", -- 3BA8
         x"c6",  x"9d",  x"cd",  x"fb",  x"b4",  x"14",  x"24",  x"e1", -- 3BB0
         x"05",  x"21",  x"03",  x"5a",  x"fb",  x"f3",  x"22",  x"e2", -- 3BB8
         x"01",  x"b5",  x"40",  x"f0",  x"3e",  x"06",  x"32",  x"cd", -- 3BC0
         x"38",  x"cd",  x"f3",  x"ae",  x"c0",  x"98",  x"fa",  x"fe", -- 3BC8
         x"54",  x"28",  x"06",  x"02",  x"fe",  x"55",  x"28",  x"1e", -- 3BD0
         x"18",  x"d8",  x"94",  x"0c",  x"6f",  x"03",  x"67",  x"a5", -- 3BD8
         x"03",  x"4f",  x"28",  x"03",  x"47",  x"03",  x"77",  x"23", -- 3BE0
         x"1f",  x"0b",  x"79",  x"b0",  x"89",  x"91",  x"18",  x"bc", -- 3BE8
         x"00",  x"1b",  x"99",  x"e1",  x"18",  x"af",  x"fb",  x"14", -- 3BF0
         x"ed",  x"4d",  x"fb",  x"70",  x"c3",  x"63",  x"b5",  x"da", -- 3BF8
         x"99",  x"9b",  x"04",  x"fe",  x"90",  x"a6",  x"04",  x"d3", -- 3C00
         x"86",  x"c2",  x"8b",  x"d3",  x"0b",  x"be",  x"58",  x"0b", -- 3C08
         x"fd",  x"b0",  x"1c",  x"ac",  x"49",  x"ec",  x"b9",  x"de", -- 3C10
         x"07",  x"8d",  x"46",  x"17",  x"e6",  x"f9",  x"1b",  x"99", -- 3C18
         x"e0",  x"18",  x"7b",  x"7c",  x"7d",  x"7e",  x"5b",  x"00", -- 3C20
         x"5c",  x"5d",  x"84",  x"94",  x"81",  x"e1",  x"8e",  x"99", -- 3C28
         x"00",  x"9a",  x"00",  x"38",  x"02",  x"03",  x"04",  x"37", -- 3C30
         x"06",  x"65",  x"07",  x"a3",  x"e0",  x"c2",  x"bd",  x"b7", -- 3C38
         x"c3",  x"69",  x"b7",  x"ce",  x"e0",  x"b3",  x"c0",  x"b7", -- 3C40
         x"c6",  x"79",  x"b7",  x"fb",  x"e0",  x"d5",  x"8e",  x"e5", -- 3C48
         x"ff",  x"68",  x"f5",  x"c5",  x"f6",  x"01",  x"f0",  x"d5", -- 3C50
         x"e3",  x"21",  x"f6",  x"77",  x"f5",  x"a6",  x"e3",  x"b1", -- 3C58
         x"86",  x"fa",  x"f1",  x"c5",  x"3a",  x"ab",  x"71",  x"da", -- 3C60
         x"e9",  x"b6",  x"92",  x"f3",  x"cf",  x"c8",  x"ce",  x"fd", -- 3C68
         x"86",  x"8f",  x"76",  x"f3",  x"b1",  x"94",  x"40",  x"f2", -- 3C70
         x"0d",  x"f2",  x"fd",  x"f1",  x"0a",  x"1a",  x"f2",  x"c7", -- 3C78
         x"f3",  x"9c",  x"e8",  x"ce",  x"4a",  x"00",  x"f7",  x"04", -- 3C80
         x"e4",  x"9b",  x"e4",  x"16",  x"e3",  x"18",  x"63",  x"e3", -- 3C88
         x"c3",  x"e7",  x"a8",  x"81",  x"20",  x"72",  x"f3",  x"5a", -- 3C90
         x"f6",  x"71",  x"00",  x"f7",  x"60",  x"f7",  x"0b",  x"f4", -- 3C98
         x"6a",  x"e0",  x"5e",  x"00",  x"e0",  x"4e",  x"e0",  x"25", -- 3CA0
         x"f9",  x"a5",  x"f4",  x"73",  x"00",  x"f8",  x"6b",  x"f8", -- 3CA8
         x"e2",  x"f6",  x"41",  x"f7",  x"41",  x"74",  x"f6",  x"91", -- 3CB0
         x"9e",  x"00",  x"f6",  x"63",  x"f8",  x"7a",  x"f7",  x"81", -- 3CB8
         x"fb",  x"79",  x"d9",  x"ad",  x"f6",  x"f7",  x"d1",  x"e9", -- 3CC0
         x"c0",  x"1c",  x"f9",  x"47",  x"f1",  x"cf",  x"62",  x"f9", -- 3CC8
         x"98",  x"57",  x"00",  x"77",  x"41",  x"61",  x"32",  x"22", -- 3CD0
         x"08",  x"19",  x"10",  x"00",  x"0c",  x"2d",  x"3d",  x"f2", -- 3CD8
         x"f8",  x"59",  x"79",  x"45",  x"01",  x"65",  x"53",  x"73", -- 3CE0
         x"33",  x"23",  x"5e",  x"5d",  x"f1",  x"ea",  x"3a",  x"2a", -- 3CE8
         x"80",  x"1d",  x"58",  x"78",  x"54",  x"74",  x"46",  x"66", -- 3CF0
         x"35",  x"00",  x"25",  x"50",  x"70",  x"1f",  x"02",  x"30", -- 3CF8
         x"40",  x"f5",  x"00",  x"fb",  x"56",  x"76",  x"55",  x"75", -- 3D00
         x"48",  x"68",  x"37",  x"01",  x"27",  x"4f",  x"6f",  x"1a", -- 3D08
         x"14",  x"39",  x"29",  x"c0",  x"ce",  x"4e",  x"6e",  x"49", -- 3D10
         x"00",  x"69",  x"4a",  x"6a",  x"38",  x"28",  x"20",  x"5b", -- 3D18
         x"4b",  x"00",  x"6b",  x"2c",  x"3c",  x"13",  x"1b",  x"4d", -- 3D20
         x"6d",  x"5a",  x"00",  x"7a",  x"47",  x"67",  x"36",  x"26", -- 3D28
         x"00",  x"00",  x"4c",  x"00",  x"6c",  x"2e",  x"3e",  x"f6", -- 3D30
         x"fc",  x"42",  x"62",  x"52",  x"00",  x"72",  x"44",  x"64", -- 3D38
         x"34",  x"24",  x"5f",  x"5c",  x"2b",  x"00",  x"3b",  x"2f", -- 3D40
         x"3f",  x"f4",  x"fa",  x"43",  x"63",  x"51",  x"00",  x"71", -- 3D48
         x"16",  x"16",  x"31",  x"21",  x"0a",  x"12",  x"0b",  x"32", -- 3D50
         x"11",  x"09",  x"cf",  x"00",  x"f7",  x"0d",  x"0d",  x"e7", -- 3D58
         x"fa",  x"08",  x"e6",  x"45",  x"62",  x"e3",  x"b5",  x"f8", -- 3D60
         x"00",  x"e5",  x"89",  x"fb",  x"39",  x"e3",  x"22",  x"e3", -- 3D68
         x"e2",  x"1c",  x"e1",  x"aa",  x"e2",  x"05",  x"a3",  x"01", -- 3D70
         x"eb",  x"e2",  x"c1",  x"0d",  x"19",  x"e1",  x"b3",  x"e1", -- 3D78
         x"90",  x"8a",  x"37",  x"e2",  x"47",  x"15",  x"07",  x"bd", -- 3D80
         x"e1",  x"45",  x"e2",  x"d6",  x"f1",  x"8d",  x"e1",  x"09", -- 3D88
         x"1a",  x"31",  x"21",  x"cb",  x"e1",  x"89",  x"17",  x"18", -- 3D90
         x"e2",  x"23",  x"06",  x"0b",  x"b1",  x"e1",  x"e5",  x"97", -- 3D98
         x"ea",  x"4e",  x"d0",  x"a1",  x"24",  x"ca",  x"4f",  x"4e", -- 3DA0
         x"f6",  x"d3",  x"6e",  x"54",  x"bf",  x"4e",  x"3f",  x"47", -- 3DA8
         x"24",  x"11",  x"0a",  x"bb",  x"f0",  x"45",  x"4e",  x"55", -- 3DB0
         x"4d",  x"6e",  x"42",  x"d0",  x"c4",  x"1c",  x"45",  x"4c", -- 3DB8
         x"45",  x"8f",  x"00",  x"d0",  x"41",  x"55",  x"53",  x"45", -- 3DC0
         x"c2",  x"45",  x"12",  x"45",  x"50",  x"d7",  x"63",  x"cb", -- 3DC8
         x"c2",  x"9e",  x"d7",  x"44",  x"1a",  x"5b",  x"39",  x"17", -- 3DD0
         x"50",  x"07",  x"17",  x"c1",  x"54",  x"c3",  x"b0",  x"ad", -- 3DD8
         x"d3",  x"86",  x"b6",  x"1b",  x"d0",  x"26",  x"54",  x"14", -- 3DE0
         x"d0",  x"52",  x"45",  x"05",  x"c2",  x"be",  x"ee",  x"66", -- 3DE8
         x"d6",  x"1e",  x"45",  x"4b",  x"04",  x"4f",  x"c3",  x"62", -- 3DF0
         x"cc",  x"4f",  x"43",  x"41",  x"47",  x"4b",  x"cb",  x"bb", -- 3DF8
         x"74",  x"06",  x"d3",  x"f4",  x"95",  x"54",  x"43",  x"3d", -- 3E00
         x"48",  x"d0",  x"12",  x"0d",  x"c3",  x"ec",  x"29",  x"2f", -- 3E08
         x"cf",  x"29",  x"4e",  x"d2",  x"50",  x"41",  x"5c",  x"4d", -- 3E10
         x"49",  x"5a",  x"19",  x"45",  x"d6",  x"47",  x"3f",  x"24", -- 3E18
         x"cc",  x"83",  x"6a",  x"45",  x"c3",  x"49",  x"52",  x"43", -- 3E20
         x"7f",  x"18",  x"c3",  x"53",  x"52",  x"35",  x"4e",  x"80", -- 3E28
         x"7d",  x"00",  x"eb",  x"fd",  x"02",  x"06",  x"e7",  x"24", -- 3E30
         x"ec",  x"65",  x"00",  x"e7",  x"45",  x"e9",  x"6a",  x"e9", -- 3E38
         x"9e",  x"e9",  x"b3",  x"00",  x"e9",  x"89",  x"ea",  x"fa", -- 3E40
         x"ea",  x"14",  x"eb",  x"48",  x"00",  x"c3",  x"30",  x"eb", -- 3E48
         x"98",  x"eb",  x"db",  x"eb",  x"0c",  x"18",  x"ec",  x"3d", -- 3E50
         x"ea",  x"0b",  x"6c",  x"ea",  x"49",  x"01",  x"eb",  x"a8", -- 3E58
         x"ec",  x"99",  x"ec",  x"ac",  x"ec",  x"81",  x"0b",  x"f8", -- 3E60
         x"ec",  x"39",  x"ed",  x"33",  x"ed",  x"87",  x"07",  x"6e", -- 3E68
         x"ed",  x"73",  x"ed",  x"de",  x"23",  x"20",  x"8f",  x"00", -- 3E70
         x"00",  x"00",  x"54",  x"80",  x"40",  x"20",  x"10",  x"08", -- 3E78
         x"04",  x"02",  x"ee",  x"e7",  x"43",  x"00",  x"81",  x"ff", -- 3E80
         x"03",  x"0b",  x"22",  x"72",  x"22",  x"3e",  x"0b",  x"00", -- 3E88
         x"12",  x"32",  x"7e",  x"32",  x"12",  x"00",  x"7e",  x"81", -- 3E90
         x"28",  x"b9",  x"a5",  x"01",  x"81",  x"55",  x"4a",  x"ff", -- 3E98
         x"01",  x"aa",  x"9b",  x"00",  x"28",  x"97",  x"01",  x"00", -- 3EA0
         x"0a",  x"3c",  x"42",  x"42",  x"7e",  x"06",  x"05",  x"10", -- 3EA8
         x"30",  x"7e",  x"30",  x"10",  x"02",  x"07",  x"08",  x"0c", -- 3EB0
         x"7e",  x"0c",  x"08",  x"f3",  x"0f",  x"00",  x"7c",  x"38", -- 3EB8
         x"10",  x"36",  x"08",  x"1c",  x"92",  x"ad",  x"00",  x"be", -- 3EC0
         x"0a",  x"30",  x"28",  x"06",  x"be",  x"58",  x"57",  x"c9", -- 3EC8
         x"28",  x"aa",  x"55",  x"43",  x"01",  x"3e",  x"7c",  x"7c", -- 3ED0
         x"3e",  x"03",  x"29",  x"f8",  x"f8",  x"1f",  x"04",  x"46", -- 3ED8
         x"00",  x"00",  x"7f",  x"30",  x"2a",  x"bf",  x"2f",  x"38", -- 3EE0
         x"00",  x"0c",  x"2a",  x"1c",  x"08",  x"7f",  x"7f",  x"9d", -- 3EE8
         x"a1",  x"0a",  x"b9",  x"85",  x"85",  x"b9",  x"66",  x"00", -- 3EF0
         x"5a",  x"5a",  x"42",  x"3c",  x"00",  x"88",  x"44",  x"22", -- 3EF8
         x"5f",  x"11",  x"03",  x"28",  x"80",  x"a7",  x"27",  x"22", -- 3F00
         x"7f",  x"05",  x"00",  x"11",  x"22",  x"44",  x"88",  x"80", -- 3F08
         x"03",  x"00",  x"01",  x"09",  x"0d",  x"7f",  x"0d",  x"09", -- 3F10
         x"c0",  x"c7",  x"90",  x"b0",  x"16",  x"fe",  x"b0",  x"90", -- 3F18
         x"87",  x"02",  x"7c",  x"06",  x"7c",  x"82",  x"46",  x"cc", -- 3F20
         x"cc",  x"33",  x"33",  x"f5",  x"03",  x"47",  x"a1",  x"12", -- 3F28
         x"00",  x"bd",  x"81",  x"82",  x"cf",  x"a5",  x"94",  x"07", -- 3F30
         x"99",  x"0f",  x"99",  x"60",  x"81",  x"a7",  x"3e",  x"16", -- 3F38
         x"60",  x"3e",  x"10",  x"c5",  x"1f",  x"0f",  x"0e",  x"e0", -- 3F40
         x"60",  x"09",  x"78",  x"0c",  x"7c",  x"cc",  x"76",  x"06", -- 3F48
         x"00",  x"e0",  x"60",  x"7c",  x"66",  x"00",  x"dc",  x"f0", -- 3F50
         x"0e",  x"0f",  x"cc",  x"c0",  x"cc",  x"78",  x"2b",  x"00", -- 3F58
         x"1c",  x"15",  x"00",  x"ec",  x"17",  x"0f",  x"fc",  x"c0", -- 3F60
         x"c1",  x"0f",  x"38",  x"6c",  x"60",  x"f0",  x"60",  x"d3", -- 3F68
         x"02",  x"0f",  x"76",  x"16",  x"19",  x"7c",  x"0c",  x"f8", -- 3F70
         x"2f",  x"6c",  x"76",  x"81",  x"2f",  x"e6",  x"00",  x"30", -- 3F78
         x"00",  x"70",  x"30",  x"8a",  x"00",  x"fc",  x"00",  x"0c", -- 3F80
         x"31",  x"6c",  x"0c",  x"19",  x"78",  x"17",  x"66",  x"6c", -- 3F88
         x"3b",  x"78",  x"6c",  x"17",  x"15",  x"ba",  x"17",  x"91", -- 3F90
         x"00",  x"fe",  x"fe",  x"d6",  x"c6",  x"a7",  x"07",  x"f8", -- 3F98
         x"1d",  x"c9",  x"00",  x"4f",  x"54",  x"26",  x"07",  x"dc", -- 3FA0
         x"dc",  x"3e",  x"7c",  x"50",  x"ca",  x"4f",  x"1e",  x"0f", -- 3FA8
         x"e4",  x"4f",  x"5f",  x"7d",  x"7c",  x"6d",  x"5e",  x"0b", -- 3FB0
         x"de",  x"7c",  x"3e",  x"2e",  x"34",  x"18",  x"3f",  x"60", -- 3FB8
         x"87",  x"bf",  x"36",  x"6d",  x"00",  x"35",  x"c6",  x"d6", -- 3FC0
         x"50",  x"6c",  x"b0",  x"07",  x"6c",  x"93",  x"be",  x"57", -- 3FC8
         x"16",  x"c3",  x"8f",  x"07",  x"0d",  x"fc",  x"98",  x"30", -- 3FD0
         x"64",  x"6f",  x"6c",  x"30",  x"cf",  x"26",  x"cc",  x"67", -- 3FD8
         x"4c",  x"cc",  x"3f",  x"3c",  x"d4",  x"6d",  x"6c",  x"02", -- 3FE0
         x"f0",  x"24",  x"ff",  x"81",  x"00",  x"40",  x"ff",  x"00", -- 3FE8
         x"20",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00", -- 3FF0
         x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00",  x"00"  -- 3FF8
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
